library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; 

entity sine_lut is 
  port (
    clk_port   : in std_logic; 
    addr       : in std_logic_vector(15 downto 0); 
    sine_out   : out std_logic_vector(15 downto 0)); -- 2.14 fixed point 
end entity sine_lut; 

architecture behavioral of sine_lut is 
  -- 2048 entries of 16 bit , 14 dec precision signed fixed point sine values 
  type rom_2048x16_t is array (0 to 2047) of std_logic_vector(15 downto 0);
  signal addr_uint : unsigned(15 downto 0) := (others => '0'); 

  -- generate table from regfile decleration 
  constant sine_table : rom_2048x16_t := (
    x"0000", x"0019", x"0032", x"004B",
    x"0065", x"007E", x"0097", x"00B0",
    x"00C9", x"00E2", x"00FB", x"0114",
    x"012E", x"0147", x"0160", x"0179",
    x"0192", x"01AB", x"01C4", x"01DD",
    x"01F7", x"0210", x"0229", x"0242",
    x"025B", x"0274", x"028D", x"02A6",
    x"02C0", x"02D9", x"02F2", x"030B",
    x"0324", x"033D", x"0356", x"036F",
    x"0388", x"03A1", x"03BB", x"03D4",
    x"03ED", x"0406", x"041F", x"0438",
    x"0451", x"046A", x"0483", x"049C",
    x"04B5", x"04CE", x"04E7", x"0500",
    x"051A", x"0533", x"054C", x"0565",
    x"057E", x"0597", x"05B0", x"05C9",
    x"05E2", x"05FB", x"0614", x"062D",
    x"0646", x"065F", x"0678", x"0691",
    x"06AA", x"06C3", x"06DC", x"06F5",
    x"070E", x"0727", x"0740", x"0759",
    x"0772", x"078B", x"07A4", x"07BD",
    x"07D6", x"07EF", x"0807", x"0820",
    x"0839", x"0852", x"086B", x"0884",
    x"089D", x"08B6", x"08CF", x"08E8",
    x"0901", x"0919", x"0932", x"094B",
    x"0964", x"097D", x"0996", x"09AF",
    x"09C7", x"09E0", x"09F9", x"0A12",
    x"0A2B", x"0A44", x"0A5C", x"0A75",
    x"0A8E", x"0AA7", x"0AC0", x"0AD8",
    x"0AF1", x"0B0A", x"0B23", x"0B3B",
    x"0B54", x"0B6D", x"0B85", x"0B9E",
    x"0BB7", x"0BD0", x"0BE8", x"0C01",
    x"0C1A", x"0C32", x"0C4B", x"0C64",
    x"0C7C", x"0C95", x"0CAE", x"0CC6",
    x"0CDF", x"0CF8", x"0D10", x"0D29",
    x"0D41", x"0D5A", x"0D72", x"0D8B",
    x"0DA4", x"0DBC", x"0DD5", x"0DED",
    x"0E06", x"0E1E", x"0E37", x"0E4F",
    x"0E68", x"0E80", x"0E99", x"0EB1",
    x"0ECA", x"0EE2", x"0EFB", x"0F13",
    x"0F2B", x"0F44", x"0F5C", x"0F75",
    x"0F8D", x"0FA5", x"0FBE", x"0FD6",
    x"0FEE", x"1007", x"101F", x"1037",
    x"1050", x"1068", x"1080", x"1099",
    x"10B1", x"10C9", x"10E1", x"10FA",
    x"1112", x"112A", x"1142", x"115A",
    x"1173", x"118B", x"11A3", x"11BB",
    x"11D3", x"11EB", x"1204", x"121C",
    x"1234", x"124C", x"1264", x"127C",
    x"1294", x"12AC", x"12C4", x"12DC",
    x"12F4", x"130C", x"1324", x"133C",
    x"1354", x"136C", x"1384", x"139C",
    x"13B4", x"13CC", x"13E4", x"13FB",
    x"1413", x"142B", x"1443", x"145B",
    x"1473", x"148B", x"14A2", x"14BA",
    x"14D2", x"14EA", x"1501", x"1519",
    x"1531", x"1549", x"1560", x"1578",
    x"1590", x"15A7", x"15BF", x"15D7",
    x"15EE", x"1606", x"161D", x"1635",
    x"164C", x"1664", x"167C", x"1693",
    x"16AB", x"16C2", x"16DA", x"16F1",
    x"1709", x"1720", x"1737", x"174F",
    x"1766", x"177E", x"1795", x"17AC",
    x"17C4", x"17DB", x"17F2", x"180A",
    x"1821", x"1838", x"184F", x"1867",
    x"187E", x"1895", x"18AC", x"18C3",
    x"18DB", x"18F2", x"1909", x"1920",
    x"1937", x"194E", x"1965", x"197C",
    x"1993", x"19AA", x"19C1", x"19D8",
    x"19EF", x"1A06", x"1A1D", x"1A34",
    x"1A4B", x"1A62", x"1A79", x"1A90",
    x"1AA7", x"1ABE", x"1AD4", x"1AEB",
    x"1B02", x"1B19", x"1B30", x"1B46",
    x"1B5D", x"1B74", x"1B8A", x"1BA1",
    x"1BB8", x"1BCE", x"1BE5", x"1BFC",
    x"1C12", x"1C29", x"1C3F", x"1C56",
    x"1C6C", x"1C83", x"1C99", x"1CB0",
    x"1CC6", x"1CDD", x"1CF3", x"1D0A",
    x"1D20", x"1D36", x"1D4D", x"1D63",
    x"1D79", x"1D90", x"1DA6", x"1DBC",
    x"1DD3", x"1DE9", x"1DFF", x"1E15",
    x"1E2B", x"1E42", x"1E58", x"1E6E",
    x"1E84", x"1E9A", x"1EB0", x"1EC6",
    x"1EDC", x"1EF2", x"1F08", x"1F1E",
    x"1F34", x"1F4A", x"1F60", x"1F76",
    x"1F8C", x"1FA2", x"1FB7", x"1FCD",
    x"1FE3", x"1FF9", x"200F", x"2024",
    x"203A", x"2050", x"2065", x"207B",
    x"2091", x"20A6", x"20BC", x"20D1",
    x"20E7", x"20FD", x"2112", x"2128",
    x"213D", x"2153", x"2168", x"217D",
    x"2193", x"21A8", x"21BE", x"21D3",
    x"21E8", x"21FE", x"2213", x"2228",
    x"223D", x"2253", x"2268", x"227D",
    x"2292", x"22A7", x"22BC", x"22D2",
    x"22E7", x"22FC", x"2311", x"2326",
    x"233B", x"2350", x"2365", x"237A",
    x"238E", x"23A3", x"23B8", x"23CD",
    x"23E2", x"23F7", x"240B", x"2420",
    x"2435", x"244A", x"245E", x"2473",
    x"2488", x"249C", x"24B1", x"24C5",
    x"24DA", x"24EF", x"2503", x"2518",
    x"252C", x"2541", x"2555", x"2569",
    x"257E", x"2592", x"25A6", x"25BB",
    x"25CF", x"25E3", x"25F8", x"260C",
    x"2620", x"2634", x"2648", x"265C",
    x"2671", x"2685", x"2699", x"26AD",
    x"26C1", x"26D5", x"26E9", x"26FD",
    x"2711", x"2724", x"2738", x"274C",
    x"2760", x"2774", x"2788", x"279B",
    x"27AF", x"27C3", x"27D6", x"27EA",
    x"27FE", x"2811", x"2825", x"2838",
    x"284C", x"2860", x"2873", x"2886",
    x"289A", x"28AD", x"28C1", x"28D4",
    x"28E7", x"28FB", x"290E", x"2921",
    x"2935", x"2948", x"295B", x"296E",
    x"2981", x"2994", x"29A7", x"29BB",
    x"29CE", x"29E1", x"29F4", x"2A07",
    x"2A1A", x"2A2C", x"2A3F", x"2A52",
    x"2A65", x"2A78", x"2A8B", x"2A9D",
    x"2AB0", x"2AC3", x"2AD6", x"2AE8",
    x"2AFB", x"2B0D", x"2B20", x"2B33",
    x"2B45", x"2B58", x"2B6A", x"2B7D",
    x"2B8F", x"2BA1", x"2BB4", x"2BC6",
    x"2BD8", x"2BEB", x"2BFD", x"2C0F",
    x"2C21", x"2C34", x"2C46", x"2C58",
    x"2C6A", x"2C7C", x"2C8E", x"2CA0",
    x"2CB2", x"2CC4", x"2CD6", x"2CE8",
    x"2CFA", x"2D0C", x"2D1E", x"2D2F",
    x"2D41", x"2D53", x"2D65", x"2D76",
    x"2D88", x"2D9A", x"2DAB", x"2DBD",
    x"2DCF", x"2DE0", x"2DF2", x"2E03",
    x"2E15", x"2E26", x"2E37", x"2E49",
    x"2E5A", x"2E6B", x"2E7D", x"2E8E",
    x"2E9F", x"2EB0", x"2EC2", x"2ED3",
    x"2EE4", x"2EF5", x"2F06", x"2F17",
    x"2F28", x"2F39", x"2F4A", x"2F5B",
    x"2F6C", x"2F7D", x"2F8D", x"2F9E",
    x"2FAF", x"2FC0", x"2FD0", x"2FE1",
    x"2FF2", x"3002", x"3013", x"3024",
    x"3034", x"3045", x"3055", x"3066",
    x"3076", x"3087", x"3097", x"30A7",
    x"30B8", x"30C8", x"30D8", x"30E8",
    x"30F9", x"3109", x"3119", x"3129",
    x"3139", x"3149", x"3159", x"3169",
    x"3179", x"3189", x"3199", x"31A9",
    x"31B9", x"31C8", x"31D8", x"31E8",
    x"31F8", x"3207", x"3217", x"3227",
    x"3236", x"3246", x"3255", x"3265",
    x"3274", x"3284", x"3293", x"32A3",
    x"32B2", x"32C1", x"32D0", x"32E0",
    x"32EF", x"32FE", x"330D", x"331D",
    x"332C", x"333B", x"334A", x"3359",
    x"3368", x"3377", x"3386", x"3395",
    x"33A3", x"33B2", x"33C1", x"33D0",
    x"33DF", x"33ED", x"33FC", x"340B",
    x"3419", x"3428", x"3436", x"3445",
    x"3453", x"3462", x"3470", x"347F",
    x"348D", x"349B", x"34AA", x"34B8",
    x"34C6", x"34D4", x"34E2", x"34F1",
    x"34FF", x"350D", x"351B", x"3529",
    x"3537", x"3545", x"3553", x"3561",
    x"356E", x"357C", x"358A", x"3598",
    x"35A5", x"35B3", x"35C1", x"35CE",
    x"35DC", x"35EA", x"35F7", x"3605",
    x"3612", x"3620", x"362D", x"363A",
    x"3648", x"3655", x"3662", x"366F",
    x"367D", x"368A", x"3697", x"36A4",
    x"36B1", x"36BE", x"36CB", x"36D8",
    x"36E5", x"36F2", x"36FF", x"370C",
    x"3718", x"3725", x"3732", x"373F",
    x"374B", x"3758", x"3765", x"3771",
    x"377E", x"378A", x"3797", x"37A3",
    x"37B0", x"37BC", x"37C8", x"37D5",
    x"37E1", x"37ED", x"37F9", x"3805",
    x"3812", x"381E", x"382A", x"3836",
    x"3842", x"384E", x"385A", x"3866",
    x"3871", x"387D", x"3889", x"3895",
    x"38A1", x"38AC", x"38B8", x"38C3",
    x"38CF", x"38DB", x"38E6", x"38F2",
    x"38FD", x"3909", x"3914", x"391F",
    x"392B", x"3936", x"3941", x"394C",
    x"3958", x"3963", x"396E", x"3979",
    x"3984", x"398F", x"399A", x"39A5",
    x"39B0", x"39BB", x"39C5", x"39D0",
    x"39DB", x"39E6", x"39F0", x"39FB",
    x"3A06", x"3A10", x"3A1B", x"3A25",
    x"3A30", x"3A3A", x"3A45", x"3A4F",
    x"3A59", x"3A64", x"3A6E", x"3A78",
    x"3A82", x"3A8D", x"3A97", x"3AA1",
    x"3AAB", x"3AB5", x"3ABF", x"3AC9",
    x"3AD3", x"3ADD", x"3AE6", x"3AF0",
    x"3AFA", x"3B04", x"3B0E", x"3B17",
    x"3B21", x"3B2A", x"3B34", x"3B3E",
    x"3B47", x"3B50", x"3B5A", x"3B63",
    x"3B6D", x"3B76", x"3B7F", x"3B88",
    x"3B92", x"3B9B", x"3BA4", x"3BAD",
    x"3BB6", x"3BBF", x"3BC8", x"3BD1",
    x"3BDA", x"3BE3", x"3BEC", x"3BF5",
    x"3BFD", x"3C06", x"3C0F", x"3C17",
    x"3C20", x"3C29", x"3C31", x"3C3A",
    x"3C42", x"3C4B", x"3C53", x"3C5B",
    x"3C64", x"3C6C", x"3C74", x"3C7D",
    x"3C85", x"3C8D", x"3C95", x"3C9D",
    x"3CA5", x"3CAD", x"3CB5", x"3CBD",
    x"3CC5", x"3CCD", x"3CD5", x"3CDD",
    x"3CE4", x"3CEC", x"3CF4", x"3CFB",
    x"3D03", x"3D0B", x"3D12", x"3D1A",
    x"3D21", x"3D28", x"3D30", x"3D37",
    x"3D3F", x"3D46", x"3D4D", x"3D54",
    x"3D5B", x"3D63", x"3D6A", x"3D71",
    x"3D78", x"3D7F", x"3D86", x"3D8D",
    x"3D93", x"3D9A", x"3DA1", x"3DA8",
    x"3DAF", x"3DB5", x"3DBC", x"3DC2",
    x"3DC9", x"3DD0", x"3DD6", x"3DDD",
    x"3DE3", x"3DE9", x"3DF0", x"3DF6",
    x"3DFC", x"3E03", x"3E09", x"3E0F",
    x"3E15", x"3E1B", x"3E21", x"3E27",
    x"3E2D", x"3E33", x"3E39", x"3E3F",
    x"3E45", x"3E4A", x"3E50", x"3E56",
    x"3E5C", x"3E61", x"3E67", x"3E6C",
    x"3E72", x"3E77", x"3E7D", x"3E82",
    x"3E88", x"3E8D", x"3E92", x"3E98",
    x"3E9D", x"3EA2", x"3EA7", x"3EAC",
    x"3EB1", x"3EB6", x"3EBB", x"3EC0",
    x"3EC5", x"3ECA", x"3ECF", x"3ED4",
    x"3ED8", x"3EDD", x"3EE2", x"3EE7",
    x"3EEB", x"3EF0", x"3EF4", x"3EF9",
    x"3EFD", x"3F02", x"3F06", x"3F0A",
    x"3F0F", x"3F13", x"3F17", x"3F1C",
    x"3F20", x"3F24", x"3F28", x"3F2C",
    x"3F30", x"3F34", x"3F38", x"3F3C",
    x"3F40", x"3F43", x"3F47", x"3F4B",
    x"3F4F", x"3F52", x"3F56", x"3F5A",
    x"3F5D", x"3F61", x"3F64", x"3F68",
    x"3F6B", x"3F6E", x"3F72", x"3F75",
    x"3F78", x"3F7B", x"3F7F", x"3F82",
    x"3F85", x"3F88", x"3F8B", x"3F8E",
    x"3F91", x"3F94", x"3F97", x"3F99",
    x"3F9C", x"3F9F", x"3FA2", x"3FA4",
    x"3FA7", x"3FAA", x"3FAC", x"3FAF",
    x"3FB1", x"3FB4", x"3FB6", x"3FB8",
    x"3FBB", x"3FBD", x"3FBF", x"3FC1",
    x"3FC4", x"3FC6", x"3FC8", x"3FCA",
    x"3FCC", x"3FCE", x"3FD0", x"3FD2",
    x"3FD4", x"3FD5", x"3FD7", x"3FD9",
    x"3FDB", x"3FDC", x"3FDE", x"3FE0",
    x"3FE1", x"3FE3", x"3FE4", x"3FE6",
    x"3FE7", x"3FE8", x"3FEA", x"3FEB",
    x"3FEC", x"3FED", x"3FEF", x"3FF0",
    x"3FF1", x"3FF2", x"3FF3", x"3FF4",
    x"3FF5", x"3FF6", x"3FF7", x"3FF7",
    x"3FF8", x"3FF9", x"3FFA", x"3FFA",
    x"3FFB", x"3FFC", x"3FFC", x"3FFD",
    x"3FFD", x"3FFE", x"3FFE", x"3FFE",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFE", x"3FFE", x"3FFE",
    x"3FFD", x"3FFD", x"3FFC", x"3FFC",
    x"3FFB", x"3FFA", x"3FFA", x"3FF9",
    x"3FF8", x"3FF7", x"3FF7", x"3FF6",
    x"3FF5", x"3FF4", x"3FF3", x"3FF2",
    x"3FF1", x"3FF0", x"3FEF", x"3FED",
    x"3FEC", x"3FEB", x"3FEA", x"3FE8",
    x"3FE7", x"3FE6", x"3FE4", x"3FE3",
    x"3FE1", x"3FE0", x"3FDE", x"3FDC",
    x"3FDB", x"3FD9", x"3FD7", x"3FD5",
    x"3FD4", x"3FD2", x"3FD0", x"3FCE",
    x"3FCC", x"3FCA", x"3FC8", x"3FC6",
    x"3FC4", x"3FC1", x"3FBF", x"3FBD",
    x"3FBB", x"3FB8", x"3FB6", x"3FB4",
    x"3FB1", x"3FAF", x"3FAC", x"3FAA",
    x"3FA7", x"3FA4", x"3FA2", x"3F9F",
    x"3F9C", x"3F99", x"3F97", x"3F94",
    x"3F91", x"3F8E", x"3F8B", x"3F88",
    x"3F85", x"3F82", x"3F7F", x"3F7B",
    x"3F78", x"3F75", x"3F72", x"3F6E",
    x"3F6B", x"3F68", x"3F64", x"3F61",
    x"3F5D", x"3F5A", x"3F56", x"3F52",
    x"3F4F", x"3F4B", x"3F47", x"3F43",
    x"3F40", x"3F3C", x"3F38", x"3F34",
    x"3F30", x"3F2C", x"3F28", x"3F24",
    x"3F20", x"3F1C", x"3F17", x"3F13",
    x"3F0F", x"3F0A", x"3F06", x"3F02",
    x"3EFD", x"3EF9", x"3EF4", x"3EF0",
    x"3EEB", x"3EE7", x"3EE2", x"3EDD",
    x"3ED8", x"3ED4", x"3ECF", x"3ECA",
    x"3EC5", x"3EC0", x"3EBB", x"3EB6",
    x"3EB1", x"3EAC", x"3EA7", x"3EA2",
    x"3E9D", x"3E98", x"3E92", x"3E8D",
    x"3E88", x"3E82", x"3E7D", x"3E77",
    x"3E72", x"3E6C", x"3E67", x"3E61",
    x"3E5C", x"3E56", x"3E50", x"3E4A",
    x"3E45", x"3E3F", x"3E39", x"3E33",
    x"3E2D", x"3E27", x"3E21", x"3E1B",
    x"3E15", x"3E0F", x"3E09", x"3E03",
    x"3DFC", x"3DF6", x"3DF0", x"3DE9",
    x"3DE3", x"3DDD", x"3DD6", x"3DD0",
    x"3DC9", x"3DC2", x"3DBC", x"3DB5",
    x"3DAF", x"3DA8", x"3DA1", x"3D9A",
    x"3D93", x"3D8D", x"3D86", x"3D7F",
    x"3D78", x"3D71", x"3D6A", x"3D63",
    x"3D5B", x"3D54", x"3D4D", x"3D46",
    x"3D3F", x"3D37", x"3D30", x"3D28",
    x"3D21", x"3D1A", x"3D12", x"3D0B",
    x"3D03", x"3CFB", x"3CF4", x"3CEC",
    x"3CE4", x"3CDD", x"3CD5", x"3CCD",
    x"3CC5", x"3CBD", x"3CB5", x"3CAD",
    x"3CA5", x"3C9D", x"3C95", x"3C8D",
    x"3C85", x"3C7D", x"3C74", x"3C6C",
    x"3C64", x"3C5B", x"3C53", x"3C4B",
    x"3C42", x"3C3A", x"3C31", x"3C29",
    x"3C20", x"3C17", x"3C0F", x"3C06",
    x"3BFD", x"3BF5", x"3BEC", x"3BE3",
    x"3BDA", x"3BD1", x"3BC8", x"3BBF",
    x"3BB6", x"3BAD", x"3BA4", x"3B9B",
    x"3B92", x"3B88", x"3B7F", x"3B76",
    x"3B6D", x"3B63", x"3B5A", x"3B50",
    x"3B47", x"3B3E", x"3B34", x"3B2A",
    x"3B21", x"3B17", x"3B0E", x"3B04",
    x"3AFA", x"3AF0", x"3AE6", x"3ADD",
    x"3AD3", x"3AC9", x"3ABF", x"3AB5",
    x"3AAB", x"3AA1", x"3A97", x"3A8D",
    x"3A82", x"3A78", x"3A6E", x"3A64",
    x"3A59", x"3A4F", x"3A45", x"3A3A",
    x"3A30", x"3A25", x"3A1B", x"3A10",
    x"3A06", x"39FB", x"39F0", x"39E6",
    x"39DB", x"39D0", x"39C5", x"39BB",
    x"39B0", x"39A5", x"399A", x"398F",
    x"3984", x"3979", x"396E", x"3963",
    x"3958", x"394C", x"3941", x"3936",
    x"392B", x"391F", x"3914", x"3909",
    x"38FD", x"38F2", x"38E6", x"38DB",
    x"38CF", x"38C3", x"38B8", x"38AC",
    x"38A1", x"3895", x"3889", x"387D",
    x"3871", x"3866", x"385A", x"384E",
    x"3842", x"3836", x"382A", x"381E",
    x"3812", x"3805", x"37F9", x"37ED",
    x"37E1", x"37D5", x"37C8", x"37BC",
    x"37B0", x"37A3", x"3797", x"378A",
    x"377E", x"3771", x"3765", x"3758",
    x"374B", x"373F", x"3732", x"3725",
    x"3718", x"370C", x"36FF", x"36F2",
    x"36E5", x"36D8", x"36CB", x"36BE",
    x"36B1", x"36A4", x"3697", x"368A",
    x"367D", x"366F", x"3662", x"3655",
    x"3648", x"363A", x"362D", x"3620",
    x"3612", x"3605", x"35F7", x"35EA",
    x"35DC", x"35CE", x"35C1", x"35B3",
    x"35A5", x"3598", x"358A", x"357C",
    x"356E", x"3561", x"3553", x"3545",
    x"3537", x"3529", x"351B", x"350D",
    x"34FF", x"34F1", x"34E2", x"34D4",
    x"34C6", x"34B8", x"34AA", x"349B",
    x"348D", x"347F", x"3470", x"3462",
    x"3453", x"3445", x"3436", x"3428",
    x"3419", x"340B", x"33FC", x"33ED",
    x"33DF", x"33D0", x"33C1", x"33B2",
    x"33A3", x"3395", x"3386", x"3377",
    x"3368", x"3359", x"334A", x"333B",
    x"332C", x"331D", x"330D", x"32FE",
    x"32EF", x"32E0", x"32D0", x"32C1",
    x"32B2", x"32A3", x"3293", x"3284",
    x"3274", x"3265", x"3255", x"3246",
    x"3236", x"3227", x"3217", x"3207",
    x"31F8", x"31E8", x"31D8", x"31C8",
    x"31B9", x"31A9", x"3199", x"3189",
    x"3179", x"3169", x"3159", x"3149",
    x"3139", x"3129", x"3119", x"3109",
    x"30F9", x"30E8", x"30D8", x"30C8",
    x"30B8", x"30A7", x"3097", x"3087",
    x"3076", x"3066", x"3055", x"3045",
    x"3034", x"3024", x"3013", x"3002",
    x"2FF2", x"2FE1", x"2FD0", x"2FC0",
    x"2FAF", x"2F9E", x"2F8D", x"2F7D",
    x"2F6C", x"2F5B", x"2F4A", x"2F39",
    x"2F28", x"2F17", x"2F06", x"2EF5",
    x"2EE4", x"2ED3", x"2EC2", x"2EB0",
    x"2E9F", x"2E8E", x"2E7D", x"2E6B",
    x"2E5A", x"2E49", x"2E37", x"2E26",
    x"2E15", x"2E03", x"2DF2", x"2DE0",
    x"2DCF", x"2DBD", x"2DAB", x"2D9A",
    x"2D88", x"2D76", x"2D65", x"2D53",
    x"2D41", x"2D2F", x"2D1E", x"2D0C",
    x"2CFA", x"2CE8", x"2CD6", x"2CC4",
    x"2CB2", x"2CA0", x"2C8E", x"2C7C",
    x"2C6A", x"2C58", x"2C46", x"2C34",
    x"2C21", x"2C0F", x"2BFD", x"2BEB",
    x"2BD8", x"2BC6", x"2BB4", x"2BA1",
    x"2B8F", x"2B7D", x"2B6A", x"2B58",
    x"2B45", x"2B33", x"2B20", x"2B0D",
    x"2AFB", x"2AE8", x"2AD6", x"2AC3",
    x"2AB0", x"2A9D", x"2A8B", x"2A78",
    x"2A65", x"2A52", x"2A3F", x"2A2C",
    x"2A1A", x"2A07", x"29F4", x"29E1",
    x"29CE", x"29BB", x"29A7", x"2994",
    x"2981", x"296E", x"295B", x"2948",
    x"2935", x"2921", x"290E", x"28FB",
    x"28E7", x"28D4", x"28C1", x"28AD",
    x"289A", x"2886", x"2873", x"2860",
    x"284C", x"2838", x"2825", x"2811",
    x"27FE", x"27EA", x"27D6", x"27C3",
    x"27AF", x"279B", x"2788", x"2774",
    x"2760", x"274C", x"2738", x"2724",
    x"2711", x"26FD", x"26E9", x"26D5",
    x"26C1", x"26AD", x"2699", x"2685",
    x"2671", x"265C", x"2648", x"2634",
    x"2620", x"260C", x"25F8", x"25E3",
    x"25CF", x"25BB", x"25A6", x"2592",
    x"257E", x"2569", x"2555", x"2541",
    x"252C", x"2518", x"2503", x"24EF",
    x"24DA", x"24C5", x"24B1", x"249C",
    x"2488", x"2473", x"245E", x"244A",
    x"2435", x"2420", x"240B", x"23F7",
    x"23E2", x"23CD", x"23B8", x"23A3",
    x"238E", x"237A", x"2365", x"2350",
    x"233B", x"2326", x"2311", x"22FC",
    x"22E7", x"22D2", x"22BC", x"22A7",
    x"2292", x"227D", x"2268", x"2253",
    x"223D", x"2228", x"2213", x"21FE",
    x"21E8", x"21D3", x"21BE", x"21A8",
    x"2193", x"217D", x"2168", x"2153",
    x"213D", x"2128", x"2112", x"20FD",
    x"20E7", x"20D1", x"20BC", x"20A6",
    x"2091", x"207B", x"2065", x"2050",
    x"203A", x"2024", x"200F", x"1FF9",
    x"1FE3", x"1FCD", x"1FB7", x"1FA2",
    x"1F8C", x"1F76", x"1F60", x"1F4A",
    x"1F34", x"1F1E", x"1F08", x"1EF2",
    x"1EDC", x"1EC6", x"1EB0", x"1E9A",
    x"1E84", x"1E6E", x"1E58", x"1E42",
    x"1E2B", x"1E15", x"1DFF", x"1DE9",
    x"1DD3", x"1DBC", x"1DA6", x"1D90",
    x"1D79", x"1D63", x"1D4D", x"1D36",
    x"1D20", x"1D0A", x"1CF3", x"1CDD",
    x"1CC6", x"1CB0", x"1C99", x"1C83",
    x"1C6C", x"1C56", x"1C3F", x"1C29",
    x"1C12", x"1BFC", x"1BE5", x"1BCE",
    x"1BB8", x"1BA1", x"1B8A", x"1B74",
    x"1B5D", x"1B46", x"1B30", x"1B19",
    x"1B02", x"1AEB", x"1AD4", x"1ABE",
    x"1AA7", x"1A90", x"1A79", x"1A62",
    x"1A4B", x"1A34", x"1A1D", x"1A06",
    x"19EF", x"19D8", x"19C1", x"19AA",
    x"1993", x"197C", x"1965", x"194E",
    x"1937", x"1920", x"1909", x"18F2",
    x"18DB", x"18C3", x"18AC", x"1895",
    x"187E", x"1867", x"184F", x"1838",
    x"1821", x"180A", x"17F2", x"17DB",
    x"17C4", x"17AC", x"1795", x"177E",
    x"1766", x"174F", x"1737", x"1720",
    x"1709", x"16F1", x"16DA", x"16C2",
    x"16AB", x"1693", x"167C", x"1664",
    x"164C", x"1635", x"161D", x"1606",
    x"15EE", x"15D7", x"15BF", x"15A7",
    x"1590", x"1578", x"1560", x"1549",
    x"1531", x"1519", x"1501", x"14EA",
    x"14D2", x"14BA", x"14A2", x"148B",
    x"1473", x"145B", x"1443", x"142B",
    x"1413", x"13FB", x"13E4", x"13CC",
    x"13B4", x"139C", x"1384", x"136C",
    x"1354", x"133C", x"1324", x"130C",
    x"12F4", x"12DC", x"12C4", x"12AC",
    x"1294", x"127C", x"1264", x"124C",
    x"1234", x"121C", x"1204", x"11EB",
    x"11D3", x"11BB", x"11A3", x"118B",
    x"1173", x"115A", x"1142", x"112A",
    x"1112", x"10FA", x"10E1", x"10C9",
    x"10B1", x"1099", x"1080", x"1068",
    x"1050", x"1037", x"101F", x"1007",
    x"0FEE", x"0FD6", x"0FBE", x"0FA5",
    x"0F8D", x"0F75", x"0F5C", x"0F44",
    x"0F2B", x"0F13", x"0EFB", x"0EE2",
    x"0ECA", x"0EB1", x"0E99", x"0E80",
    x"0E68", x"0E4F", x"0E37", x"0E1E",
    x"0E06", x"0DED", x"0DD5", x"0DBC",
    x"0DA4", x"0D8B", x"0D72", x"0D5A",
    x"0D41", x"0D29", x"0D10", x"0CF8",
    x"0CDF", x"0CC6", x"0CAE", x"0C95",
    x"0C7C", x"0C64", x"0C4B", x"0C32",
    x"0C1A", x"0C01", x"0BE8", x"0BD0",
    x"0BB7", x"0B9E", x"0B85", x"0B6D",
    x"0B54", x"0B3B", x"0B23", x"0B0A",
    x"0AF1", x"0AD8", x"0AC0", x"0AA7",
    x"0A8E", x"0A75", x"0A5C", x"0A44",
    x"0A2B", x"0A12", x"09F9", x"09E0",
    x"09C7", x"09AF", x"0996", x"097D",
    x"0964", x"094B", x"0932", x"0919",
    x"0901", x"08E8", x"08CF", x"08B6",
    x"089D", x"0884", x"086B", x"0852",
    x"0839", x"0820", x"0807", x"07EF",
    x"07D6", x"07BD", x"07A4", x"078B",
    x"0772", x"0759", x"0740", x"0727",
    x"070E", x"06F5", x"06DC", x"06C3",
    x"06AA", x"0691", x"0678", x"065F",
    x"0646", x"062D", x"0614", x"05FB",
    x"05E2", x"05C9", x"05B0", x"0597",
    x"057E", x"0565", x"054C", x"0533",
    x"051A", x"0500", x"04E7", x"04CE",
    x"04B5", x"049C", x"0483", x"046A",
    x"0451", x"0438", x"041F", x"0406",
    x"03ED", x"03D4", x"03BB", x"03A1",
    x"0388", x"036F", x"0356", x"033D",
    x"0324", x"030B", x"02F2", x"02D9",
    x"02C0", x"02A6", x"028D", x"0274",
    x"025B", x"0242", x"0229", x"0210",
    x"01F7", x"01DD", x"01C4", x"01AB",
    x"0192", x"0179", x"0160", x"0147",
    x"012E", x"0114", x"00FB", x"00E2",
    x"00C9", x"00B0", x"0097", x"007E",
    x"0065", x"004B", x"0032", x"0019",
    x"0000", x"FFE7", x"FFCE", x"FFB5",
    x"FF9B", x"FF82", x"FF69", x"FF50",
    x"FF37", x"FF1E", x"FF05", x"FEEC",
    x"FED2", x"FEB9", x"FEA0", x"FE87",
    x"FE6E", x"FE55", x"FE3C", x"FE23",
    x"FE09", x"FDF0", x"FDD7", x"FDBE",
    x"FDA5", x"FD8C", x"FD73", x"FD5A",
    x"FD40", x"FD27", x"FD0E", x"FCF5",
    x"FCDC", x"FCC3", x"FCAA", x"FC91",
    x"FC78", x"FC5F", x"FC45", x"FC2C",
    x"FC13", x"FBFA", x"FBE1", x"FBC8",
    x"FBAF", x"FB96", x"FB7D", x"FB64",
    x"FB4B", x"FB32", x"FB19", x"FB00",
    x"FAE6", x"FACD", x"FAB4", x"FA9B",
    x"FA82", x"FA69", x"FA50", x"FA37",
    x"FA1E", x"FA05", x"F9EC", x"F9D3",
    x"F9BA", x"F9A1", x"F988", x"F96F",
    x"F956", x"F93D", x"F924", x"F90B",
    x"F8F2", x"F8D9", x"F8C0", x"F8A7",
    x"F88E", x"F875", x"F85C", x"F843",
    x"F82A", x"F811", x"F7F9", x"F7E0",
    x"F7C7", x"F7AE", x"F795", x"F77C",
    x"F763", x"F74A", x"F731", x"F718",
    x"F6FF", x"F6E7", x"F6CE", x"F6B5",
    x"F69C", x"F683", x"F66A", x"F651",
    x"F639", x"F620", x"F607", x"F5EE",
    x"F5D5", x"F5BC", x"F5A4", x"F58B",
    x"F572", x"F559", x"F540", x"F528",
    x"F50F", x"F4F6", x"F4DD", x"F4C5",
    x"F4AC", x"F493", x"F47B", x"F462",
    x"F449", x"F430", x"F418", x"F3FF",
    x"F3E6", x"F3CE", x"F3B5", x"F39C",
    x"F384", x"F36B", x"F352", x"F33A",
    x"F321", x"F308", x"F2F0", x"F2D7",
    x"F2BF", x"F2A6", x"F28E", x"F275",
    x"F25C", x"F244", x"F22B", x"F213",
    x"F1FA", x"F1E2", x"F1C9", x"F1B1",
    x"F198", x"F180", x"F167", x"F14F",
    x"F136", x"F11E", x"F105", x"F0ED",
    x"F0D5", x"F0BC", x"F0A4", x"F08B",
    x"F073", x"F05B", x"F042", x"F02A",
    x"F012", x"EFF9", x"EFE1", x"EFC9",
    x"EFB0", x"EF98", x"EF80", x"EF67",
    x"EF4F", x"EF37", x"EF1F", x"EF06",
    x"EEEE", x"EED6", x"EEBE", x"EEA6",
    x"EE8D", x"EE75", x"EE5D", x"EE45",
    x"EE2D", x"EE15", x"EDFC", x"EDE4",
    x"EDCC", x"EDB4", x"ED9C", x"ED84",
    x"ED6C", x"ED54", x"ED3C", x"ED24",
    x"ED0C", x"ECF4", x"ECDC", x"ECC4",
    x"ECAC", x"EC94", x"EC7C", x"EC64",
    x"EC4C", x"EC34", x"EC1C", x"EC05",
    x"EBED", x"EBD5", x"EBBD", x"EBA5",
    x"EB8D", x"EB75", x"EB5E", x"EB46",
    x"EB2E", x"EB16", x"EAFF", x"EAE7",
    x"EACF", x"EAB7", x"EAA0", x"EA88",
    x"EA70", x"EA59", x"EA41", x"EA29",
    x"EA12", x"E9FA", x"E9E3", x"E9CB",
    x"E9B4", x"E99C", x"E984", x"E96D",
    x"E955", x"E93E", x"E926", x"E90F",
    x"E8F7", x"E8E0", x"E8C9", x"E8B1",
    x"E89A", x"E882", x"E86B", x"E854",
    x"E83C", x"E825", x"E80E", x"E7F6",
    x"E7DF", x"E7C8", x"E7B1", x"E799",
    x"E782", x"E76B", x"E754", x"E73D",
    x"E725", x"E70E", x"E6F7", x"E6E0",
    x"E6C9", x"E6B2", x"E69B", x"E684",
    x"E66D", x"E656", x"E63F", x"E628",
    x"E611", x"E5FA", x"E5E3", x"E5CC",
    x"E5B5", x"E59E", x"E587", x"E570",
    x"E559", x"E542", x"E52C", x"E515",
    x"E4FE", x"E4E7", x"E4D0", x"E4BA",
    x"E4A3", x"E48C", x"E476", x"E45F",
    x"E448", x"E432", x"E41B", x"E404",
    x"E3EE", x"E3D7", x"E3C1", x"E3AA",
    x"E394", x"E37D", x"E367", x"E350",
    x"E33A", x"E323", x"E30D", x"E2F6",
    x"E2E0", x"E2CA", x"E2B3", x"E29D",
    x"E287", x"E270", x"E25A", x"E244",
    x"E22D", x"E217", x"E201", x"E1EB",
    x"E1D5", x"E1BE", x"E1A8", x"E192",
    x"E17C", x"E166", x"E150", x"E13A",
    x"E124", x"E10E", x"E0F8", x"E0E2",
    x"E0CC", x"E0B6", x"E0A0", x"E08A",
    x"E074", x"E05E", x"E049", x"E033",
    x"E01D", x"E007", x"DFF1", x"DFDC",
    x"DFC6", x"DFB0", x"DF9B", x"DF85",
    x"DF6F", x"DF5A", x"DF44", x"DF2F",
    x"DF19", x"DF03", x"DEEE", x"DED8",
    x"DEC3", x"DEAD", x"DE98", x"DE83",
    x"DE6D", x"DE58", x"DE42", x"DE2D",
    x"DE18", x"DE02", x"DDED", x"DDD8",
    x"DDC3", x"DDAD", x"DD98", x"DD83",
    x"DD6E", x"DD59", x"DD44", x"DD2E",
    x"DD19", x"DD04", x"DCEF", x"DCDA",
    x"DCC5", x"DCB0", x"DC9B", x"DC86",
    x"DC72", x"DC5D", x"DC48", x"DC33",
    x"DC1E", x"DC09", x"DBF5", x"DBE0",
    x"DBCB", x"DBB6", x"DBA2", x"DB8D",
    x"DB78", x"DB64", x"DB4F", x"DB3B",
    x"DB26", x"DB11", x"DAFD", x"DAE8",
    x"DAD4", x"DABF", x"DAAB", x"DA97",
    x"DA82", x"DA6E", x"DA5A", x"DA45",
    x"DA31", x"DA1D", x"DA08", x"D9F4",
    x"D9E0", x"D9CC", x"D9B8", x"D9A4",
    x"D98F", x"D97B", x"D967", x"D953",
    x"D93F", x"D92B", x"D917", x"D903",
    x"D8EF", x"D8DC", x"D8C8", x"D8B4",
    x"D8A0", x"D88C", x"D878", x"D865",
    x"D851", x"D83D", x"D82A", x"D816",
    x"D802", x"D7EF", x"D7DB", x"D7C8",
    x"D7B4", x"D7A0", x"D78D", x"D77A",
    x"D766", x"D753", x"D73F", x"D72C",
    x"D719", x"D705", x"D6F2", x"D6DF",
    x"D6CB", x"D6B8", x"D6A5", x"D692",
    x"D67F", x"D66C", x"D659", x"D645",
    x"D632", x"D61F", x"D60C", x"D5F9",
    x"D5E6", x"D5D4", x"D5C1", x"D5AE",
    x"D59B", x"D588", x"D575", x"D563",
    x"D550", x"D53D", x"D52A", x"D518",
    x"D505", x"D4F3", x"D4E0", x"D4CD",
    x"D4BB", x"D4A8", x"D496", x"D483",
    x"D471", x"D45F", x"D44C", x"D43A",
    x"D428", x"D415", x"D403", x"D3F1",
    x"D3DF", x"D3CC", x"D3BA", x"D3A8",
    x"D396", x"D384", x"D372", x"D360",
    x"D34E", x"D33C", x"D32A", x"D318",
    x"D306", x"D2F4", x"D2E2", x"D2D1",
    x"D2BF", x"D2AD", x"D29B", x"D28A",
    x"D278", x"D266", x"D255", x"D243",
    x"D231", x"D220", x"D20E", x"D1FD",
    x"D1EB", x"D1DA", x"D1C9", x"D1B7",
    x"D1A6", x"D195", x"D183", x"D172",
    x"D161", x"D150", x"D13E", x"D12D",
    x"D11C", x"D10B", x"D0FA", x"D0E9",
    x"D0D8", x"D0C7", x"D0B6", x"D0A5",
    x"D094", x"D083", x"D073", x"D062",
    x"D051", x"D040", x"D030", x"D01F",
    x"D00E", x"CFFE", x"CFED", x"CFDC",
    x"CFCC", x"CFBB", x"CFAB", x"CF9A",
    x"CF8A", x"CF79", x"CF69", x"CF59",
    x"CF48", x"CF38", x"CF28", x"CF18",
    x"CF07", x"CEF7", x"CEE7", x"CED7",
    x"CEC7", x"CEB7", x"CEA7", x"CE97",
    x"CE87", x"CE77", x"CE67", x"CE57",
    x"CE47", x"CE38", x"CE28", x"CE18",
    x"CE08", x"CDF9", x"CDE9", x"CDD9",
    x"CDCA", x"CDBA", x"CDAB", x"CD9B",
    x"CD8C", x"CD7C", x"CD6D", x"CD5D",
    x"CD4E", x"CD3F", x"CD30", x"CD20",
    x"CD11", x"CD02", x"CCF3", x"CCE3",
    x"CCD4", x"CCC5", x"CCB6", x"CCA7",
    x"CC98", x"CC89", x"CC7A", x"CC6B",
    x"CC5D", x"CC4E", x"CC3F", x"CC30",
    x"CC21", x"CC13", x"CC04", x"CBF5",
    x"CBE7", x"CBD8", x"CBCA", x"CBBB",
    x"CBAD", x"CB9E", x"CB90", x"CB81",
    x"CB73", x"CB65", x"CB56", x"CB48",
    x"CB3A", x"CB2C", x"CB1E", x"CB0F",
    x"CB01", x"CAF3", x"CAE5", x"CAD7",
    x"CAC9", x"CABB", x"CAAD", x"CA9F",
    x"CA92", x"CA84", x"CA76", x"CA68",
    x"CA5B", x"CA4D", x"CA3F", x"CA32",
    x"CA24", x"CA16", x"CA09", x"C9FB",
    x"C9EE", x"C9E0", x"C9D3", x"C9C6",
    x"C9B8", x"C9AB", x"C99E", x"C991",
    x"C983", x"C976", x"C969", x"C95C",
    x"C94F", x"C942", x"C935", x"C928",
    x"C91B", x"C90E", x"C901", x"C8F4",
    x"C8E8", x"C8DB", x"C8CE", x"C8C1",
    x"C8B5", x"C8A8", x"C89B", x"C88F",
    x"C882", x"C876", x"C869", x"C85D",
    x"C850", x"C844", x"C838", x"C82B",
    x"C81F", x"C813", x"C807", x"C7FB",
    x"C7EE", x"C7E2", x"C7D6", x"C7CA",
    x"C7BE", x"C7B2", x"C7A6", x"C79A",
    x"C78F", x"C783", x"C777", x"C76B",
    x"C75F", x"C754", x"C748", x"C73D",
    x"C731", x"C725", x"C71A", x"C70E",
    x"C703", x"C6F7", x"C6EC", x"C6E1",
    x"C6D5", x"C6CA", x"C6BF", x"C6B4",
    x"C6A8", x"C69D", x"C692", x"C687",
    x"C67C", x"C671", x"C666", x"C65B",
    x"C650", x"C645", x"C63B", x"C630",
    x"C625", x"C61A", x"C610", x"C605",
    x"C5FA", x"C5F0", x"C5E5", x"C5DB",
    x"C5D0", x"C5C6", x"C5BB", x"C5B1",
    x"C5A7", x"C59C", x"C592", x"C588",
    x"C57E", x"C573", x"C569", x"C55F",
    x"C555", x"C54B", x"C541", x"C537",
    x"C52D", x"C523", x"C51A", x"C510",
    x"C506", x"C4FC", x"C4F2", x"C4E9",
    x"C4DF", x"C4D6", x"C4CC", x"C4C2",
    x"C4B9", x"C4B0", x"C4A6", x"C49D",
    x"C493", x"C48A", x"C481", x"C478",
    x"C46E", x"C465", x"C45C", x"C453",
    x"C44A", x"C441", x"C438", x"C42F",
    x"C426", x"C41D", x"C414", x"C40B",
    x"C403", x"C3FA", x"C3F1", x"C3E9",
    x"C3E0", x"C3D7", x"C3CF", x"C3C6",
    x"C3BE", x"C3B5", x"C3AD", x"C3A5",
    x"C39C", x"C394", x"C38C", x"C383",
    x"C37B", x"C373", x"C36B", x"C363",
    x"C35B", x"C353", x"C34B", x"C343",
    x"C33B", x"C333", x"C32B", x"C323",
    x"C31C", x"C314", x"C30C", x"C305",
    x"C2FD", x"C2F5", x"C2EE", x"C2E6",
    x"C2DF", x"C2D8", x"C2D0", x"C2C9",
    x"C2C1", x"C2BA", x"C2B3", x"C2AC",
    x"C2A5", x"C29D", x"C296", x"C28F",
    x"C288", x"C281", x"C27A", x"C273",
    x"C26D", x"C266", x"C25F", x"C258",
    x"C251", x"C24B", x"C244", x"C23E",
    x"C237", x"C230", x"C22A", x"C223",
    x"C21D", x"C217", x"C210", x"C20A",
    x"C204", x"C1FD", x"C1F7", x"C1F1",
    x"C1EB", x"C1E5", x"C1DF", x"C1D9",
    x"C1D3", x"C1CD", x"C1C7", x"C1C1",
    x"C1BB", x"C1B6", x"C1B0", x"C1AA",
    x"C1A4", x"C19F", x"C199", x"C194",
    x"C18E", x"C189", x"C183", x"C17E",
    x"C178", x"C173", x"C16E", x"C168",
    x"C163", x"C15E", x"C159", x"C154",
    x"C14F", x"C14A", x"C145", x"C140",
    x"C13B", x"C136", x"C131", x"C12C",
    x"C128", x"C123", x"C11E", x"C119",
    x"C115", x"C110", x"C10C", x"C107",
    x"C103", x"C0FE", x"C0FA", x"C0F6",
    x"C0F1", x"C0ED", x"C0E9", x"C0E4",
    x"C0E0", x"C0DC", x"C0D8", x"C0D4",
    x"C0D0", x"C0CC", x"C0C8", x"C0C4",
    x"C0C0", x"C0BD", x"C0B9", x"C0B5",
    x"C0B1", x"C0AE", x"C0AA", x"C0A6",
    x"C0A3", x"C09F", x"C09C", x"C098",
    x"C095", x"C092", x"C08E", x"C08B",
    x"C088", x"C085", x"C081", x"C07E",
    x"C07B", x"C078", x"C075", x"C072",
    x"C06F", x"C06C", x"C069", x"C067",
    x"C064", x"C061", x"C05E", x"C05C",
    x"C059", x"C056", x"C054", x"C051",
    x"C04F", x"C04C", x"C04A", x"C048",
    x"C045", x"C043", x"C041", x"C03F",
    x"C03C", x"C03A", x"C038", x"C036",
    x"C034", x"C032", x"C030", x"C02E",
    x"C02C", x"C02B", x"C029", x"C027",
    x"C025", x"C024", x"C022", x"C020",
    x"C01F", x"C01D", x"C01C", x"C01A",
    x"C019", x"C018", x"C016", x"C015",
    x"C014", x"C013", x"C011", x"C010",
    x"C00F", x"C00E", x"C00D", x"C00C",
    x"C00B", x"C00A", x"C009", x"C009",
    x"C008", x"C007", x"C006", x"C006",
    x"C005", x"C004", x"C004", x"C003",
    x"C003", x"C002", x"C002", x"C002",
    x"C001", x"C001", x"C001", x"C000",
    x"C000", x"C000", x"C000", x"C000",
    x"C000", x"C000", x"C000", x"C000",
    x"C000", x"C000", x"C001", x"C001",
    x"C001", x"C002", x"C002", x"C002",
    x"C003", x"C003", x"C004", x"C004",
    x"C005", x"C006", x"C006", x"C007",
    x"C008", x"C009", x"C009", x"C00A",
    x"C00B", x"C00C", x"C00D", x"C00E",
    x"C00F", x"C010", x"C011", x"C013",
    x"C014", x"C015", x"C016", x"C018",
    x"C019", x"C01A", x"C01C", x"C01D",
    x"C01F", x"C020", x"C022", x"C024",
    x"C025", x"C027", x"C029", x"C02B",
    x"C02C", x"C02E", x"C030", x"C032",
    x"C034", x"C036", x"C038", x"C03A",
    x"C03C", x"C03F", x"C041", x"C043",
    x"C045", x"C048", x"C04A", x"C04C",
    x"C04F", x"C051", x"C054", x"C056",
    x"C059", x"C05C", x"C05E", x"C061",
    x"C064", x"C067", x"C069", x"C06C",
    x"C06F", x"C072", x"C075", x"C078",
    x"C07B", x"C07E", x"C081", x"C085",
    x"C088", x"C08B", x"C08E", x"C092",
    x"C095", x"C098", x"C09C", x"C09F",
    x"C0A3", x"C0A6", x"C0AA", x"C0AE",
    x"C0B1", x"C0B5", x"C0B9", x"C0BD",
    x"C0C0", x"C0C4", x"C0C8", x"C0CC",
    x"C0D0", x"C0D4", x"C0D8", x"C0DC",
    x"C0E0", x"C0E4", x"C0E9", x"C0ED",
    x"C0F1", x"C0F6", x"C0FA", x"C0FE",
    x"C103", x"C107", x"C10C", x"C110",
    x"C115", x"C119", x"C11E", x"C123",
    x"C128", x"C12C", x"C131", x"C136",
    x"C13B", x"C140", x"C145", x"C14A",
    x"C14F", x"C154", x"C159", x"C15E",
    x"C163", x"C168", x"C16E", x"C173",
    x"C178", x"C17E", x"C183", x"C189",
    x"C18E", x"C194", x"C199", x"C19F",
    x"C1A4", x"C1AA", x"C1B0", x"C1B6",
    x"C1BB", x"C1C1", x"C1C7", x"C1CD",
    x"C1D3", x"C1D9", x"C1DF", x"C1E5",
    x"C1EB", x"C1F1", x"C1F7", x"C1FD",
    x"C204", x"C20A", x"C210", x"C217",
    x"C21D", x"C223", x"C22A", x"C230",
    x"C237", x"C23E", x"C244", x"C24B",
    x"C251", x"C258", x"C25F", x"C266",
    x"C26D", x"C273", x"C27A", x"C281",
    x"C288", x"C28F", x"C296", x"C29D",
    x"C2A5", x"C2AC", x"C2B3", x"C2BA",
    x"C2C1", x"C2C9", x"C2D0", x"C2D8",
    x"C2DF", x"C2E6", x"C2EE", x"C2F5",
    x"C2FD", x"C305", x"C30C", x"C314",
    x"C31C", x"C323", x"C32B", x"C333",
    x"C33B", x"C343", x"C34B", x"C353",
    x"C35B", x"C363", x"C36B", x"C373",
    x"C37B", x"C383", x"C38C", x"C394",
    x"C39C", x"C3A5", x"C3AD", x"C3B5",
    x"C3BE", x"C3C6", x"C3CF", x"C3D7",
    x"C3E0", x"C3E9", x"C3F1", x"C3FA",
    x"C403", x"C40B", x"C414", x"C41D",
    x"C426", x"C42F", x"C438", x"C441",
    x"C44A", x"C453", x"C45C", x"C465",
    x"C46E", x"C478", x"C481", x"C48A",
    x"C493", x"C49D", x"C4A6", x"C4B0",
    x"C4B9", x"C4C2", x"C4CC", x"C4D6",
    x"C4DF", x"C4E9", x"C4F2", x"C4FC",
    x"C506", x"C510", x"C51A", x"C523",
    x"C52D", x"C537", x"C541", x"C54B",
    x"C555", x"C55F", x"C569", x"C573",
    x"C57E", x"C588", x"C592", x"C59C",
    x"C5A7", x"C5B1", x"C5BB", x"C5C6",
    x"C5D0", x"C5DB", x"C5E5", x"C5F0",
    x"C5FA", x"C605", x"C610", x"C61A",
    x"C625", x"C630", x"C63B", x"C645",
    x"C650", x"C65B", x"C666", x"C671",
    x"C67C", x"C687", x"C692", x"C69D",
    x"C6A8", x"C6B4", x"C6BF", x"C6CA",
    x"C6D5", x"C6E1", x"C6EC", x"C6F7",
    x"C703", x"C70E", x"C71A", x"C725",
    x"C731", x"C73D", x"C748", x"C754",
    x"C75F", x"C76B", x"C777", x"C783",
    x"C78F", x"C79A", x"C7A6", x"C7B2",
    x"C7BE", x"C7CA", x"C7D6", x"C7E2",
    x"C7EE", x"C7FB", x"C807", x"C813",
    x"C81F", x"C82B", x"C838", x"C844",
    x"C850", x"C85D", x"C869", x"C876",
    x"C882", x"C88F", x"C89B", x"C8A8",
    x"C8B5", x"C8C1", x"C8CE", x"C8DB",
    x"C8E8", x"C8F4", x"C901", x"C90E",
    x"C91B", x"C928", x"C935", x"C942",
    x"C94F", x"C95C", x"C969", x"C976",
    x"C983", x"C991", x"C99E", x"C9AB",
    x"C9B8", x"C9C6", x"C9D3", x"C9E0",
    x"C9EE", x"C9FB", x"CA09", x"CA16",
    x"CA24", x"CA32", x"CA3F", x"CA4D",
    x"CA5B", x"CA68", x"CA76", x"CA84",
    x"CA92", x"CA9F", x"CAAD", x"CABB",
    x"CAC9", x"CAD7", x"CAE5", x"CAF3",
    x"CB01", x"CB0F", x"CB1E", x"CB2C",
    x"CB3A", x"CB48", x"CB56", x"CB65",
    x"CB73", x"CB81", x"CB90", x"CB9E",
    x"CBAD", x"CBBB", x"CBCA", x"CBD8",
    x"CBE7", x"CBF5", x"CC04", x"CC13",
    x"CC21", x"CC30", x"CC3F", x"CC4E",
    x"CC5D", x"CC6B", x"CC7A", x"CC89",
    x"CC98", x"CCA7", x"CCB6", x"CCC5",
    x"CCD4", x"CCE3", x"CCF3", x"CD02",
    x"CD11", x"CD20", x"CD30", x"CD3F",
    x"CD4E", x"CD5D", x"CD6D", x"CD7C",
    x"CD8C", x"CD9B", x"CDAB", x"CDBA",
    x"CDCA", x"CDD9", x"CDE9", x"CDF9",
    x"CE08", x"CE18", x"CE28", x"CE38",
    x"CE47", x"CE57", x"CE67", x"CE77",
    x"CE87", x"CE97", x"CEA7", x"CEB7",
    x"CEC7", x"CED7", x"CEE7", x"CEF7",
    x"CF07", x"CF18", x"CF28", x"CF38",
    x"CF48", x"CF59", x"CF69", x"CF79",
    x"CF8A", x"CF9A", x"CFAB", x"CFBB",
    x"CFCC", x"CFDC", x"CFED", x"CFFE",
    x"D00E", x"D01F", x"D030", x"D040",
    x"D051", x"D062", x"D073", x"D083",
    x"D094", x"D0A5", x"D0B6", x"D0C7",
    x"D0D8", x"D0E9", x"D0FA", x"D10B",
    x"D11C", x"D12D", x"D13E", x"D150",
    x"D161", x"D172", x"D183", x"D195",
    x"D1A6", x"D1B7", x"D1C9", x"D1DA",
    x"D1EB", x"D1FD", x"D20E", x"D220",
    x"D231", x"D243", x"D255", x"D266",
    x"D278", x"D28A", x"D29B", x"D2AD",
    x"D2BF", x"D2D1", x"D2E2", x"D2F4",
    x"D306", x"D318", x"D32A", x"D33C",
    x"D34E", x"D360", x"D372", x"D384",
    x"D396", x"D3A8", x"D3BA", x"D3CC",
    x"D3DF", x"D3F1", x"D403", x"D415",
    x"D428", x"D43A", x"D44C", x"D45F",
    x"D471", x"D483", x"D496", x"D4A8",
    x"D4BB", x"D4CD", x"D4E0", x"D4F3",
    x"D505", x"D518", x"D52A", x"D53D",
    x"D550", x"D563", x"D575", x"D588",
    x"D59B", x"D5AE", x"D5C1", x"D5D4",
    x"D5E6", x"D5F9", x"D60C", x"D61F",
    x"D632", x"D645", x"D659", x"D66C",
    x"D67F", x"D692", x"D6A5", x"D6B8",
    x"D6CB", x"D6DF", x"D6F2", x"D705",
    x"D719", x"D72C", x"D73F", x"D753",
    x"D766", x"D77A", x"D78D", x"D7A0",
    x"D7B4", x"D7C8", x"D7DB", x"D7EF",
    x"D802", x"D816", x"D82A", x"D83D",
    x"D851", x"D865", x"D878", x"D88C",
    x"D8A0", x"D8B4", x"D8C8", x"D8DC",
    x"D8EF", x"D903", x"D917", x"D92B",
    x"D93F", x"D953", x"D967", x"D97B",
    x"D98F", x"D9A4", x"D9B8", x"D9CC",
    x"D9E0", x"D9F4", x"DA08", x"DA1D",
    x"DA31", x"DA45", x"DA5A", x"DA6E",
    x"DA82", x"DA97", x"DAAB", x"DABF",
    x"DAD4", x"DAE8", x"DAFD", x"DB11",
    x"DB26", x"DB3B", x"DB4F", x"DB64",
    x"DB78", x"DB8D", x"DBA2", x"DBB6",
    x"DBCB", x"DBE0", x"DBF5", x"DC09",
    x"DC1E", x"DC33", x"DC48", x"DC5D",
    x"DC72", x"DC86", x"DC9B", x"DCB0",
    x"DCC5", x"DCDA", x"DCEF", x"DD04",
    x"DD19", x"DD2E", x"DD44", x"DD59",
    x"DD6E", x"DD83", x"DD98", x"DDAD",
    x"DDC3", x"DDD8", x"DDED", x"DE02",
    x"DE18", x"DE2D", x"DE42", x"DE58",
    x"DE6D", x"DE83", x"DE98", x"DEAD",
    x"DEC3", x"DED8", x"DEEE", x"DF03",
    x"DF19", x"DF2F", x"DF44", x"DF5A",
    x"DF6F", x"DF85", x"DF9B", x"DFB0",
    x"DFC6", x"DFDC", x"DFF1", x"E007",
    x"E01D", x"E033", x"E049", x"E05E",
    x"E074", x"E08A", x"E0A0", x"E0B6",
    x"E0CC", x"E0E2", x"E0F8", x"E10E",
    x"E124", x"E13A", x"E150", x"E166",
    x"E17C", x"E192", x"E1A8", x"E1BE",
    x"E1D5", x"E1EB", x"E201", x"E217",
    x"E22D", x"E244", x"E25A", x"E270",
    x"E287", x"E29D", x"E2B3", x"E2CA",
    x"E2E0", x"E2F6", x"E30D", x"E323",
    x"E33A", x"E350", x"E367", x"E37D",
    x"E394", x"E3AA", x"E3C1", x"E3D7",
    x"E3EE", x"E404", x"E41B", x"E432",
    x"E448", x"E45F", x"E476", x"E48C",
    x"E4A3", x"E4BA", x"E4D0", x"E4E7",
    x"E4FE", x"E515", x"E52C", x"E542",
    x"E559", x"E570", x"E587", x"E59E",
    x"E5B5", x"E5CC", x"E5E3", x"E5FA",
    x"E611", x"E628", x"E63F", x"E656",
    x"E66D", x"E684", x"E69B", x"E6B2",
    x"E6C9", x"E6E0", x"E6F7", x"E70E",
    x"E725", x"E73D", x"E754", x"E76B",
    x"E782", x"E799", x"E7B1", x"E7C8",
    x"E7DF", x"E7F6", x"E80E", x"E825",
    x"E83C", x"E854", x"E86B", x"E882",
    x"E89A", x"E8B1", x"E8C9", x"E8E0",
    x"E8F7", x"E90F", x"E926", x"E93E",
    x"E955", x"E96D", x"E984", x"E99C",
    x"E9B4", x"E9CB", x"E9E3", x"E9FA",
    x"EA12", x"EA29", x"EA41", x"EA59",
    x"EA70", x"EA88", x"EAA0", x"EAB7",
    x"EACF", x"EAE7", x"EAFF", x"EB16",
    x"EB2E", x"EB46", x"EB5E", x"EB75",
    x"EB8D", x"EBA5", x"EBBD", x"EBD5",
    x"EBED", x"EC05", x"EC1C", x"EC34",
    x"EC4C", x"EC64", x"EC7C", x"EC94",
    x"ECAC", x"ECC4", x"ECDC", x"ECF4",
    x"ED0C", x"ED24", x"ED3C", x"ED54",
    x"ED6C", x"ED84", x"ED9C", x"EDB4",
    x"EDCC", x"EDE4", x"EDFC", x"EE15",
    x"EE2D", x"EE45", x"EE5D", x"EE75",
    x"EE8D", x"EEA6", x"EEBE", x"EED6",
    x"EEEE", x"EF06", x"EF1F", x"EF37",
    x"EF4F", x"EF67", x"EF80", x"EF98",
    x"EFB0", x"EFC9", x"EFE1", x"EFF9",
    x"F012", x"F02A", x"F042", x"F05B",
    x"F073", x"F08B", x"F0A4", x"F0BC",
    x"F0D5", x"F0ED", x"F105", x"F11E",
    x"F136", x"F14F", x"F167", x"F180",
    x"F198", x"F1B1", x"F1C9", x"F1E2",
    x"F1FA", x"F213", x"F22B", x"F244",
    x"F25C", x"F275", x"F28E", x"F2A6",
    x"F2BF", x"F2D7", x"F2F0", x"F308",
    x"F321", x"F33A", x"F352", x"F36B",
    x"F384", x"F39C", x"F3B5", x"F3CE",
    x"F3E6", x"F3FF", x"F418", x"F430",
    x"F449", x"F462", x"F47B", x"F493",
    x"F4AC", x"F4C5", x"F4DD", x"F4F6",
    x"F50F", x"F528", x"F540", x"F559",
    x"F572", x"F58B", x"F5A4", x"F5BC",
    x"F5D5", x"F5EE", x"F607", x"F620",
    x"F639", x"F651", x"F66A", x"F683",
    x"F69C", x"F6B5", x"F6CE", x"F6E7",
    x"F6FF", x"F718", x"F731", x"F74A",
    x"F763", x"F77C", x"F795", x"F7AE",
    x"F7C7", x"F7E0", x"F7F9", x"F811",
    x"F82A", x"F843", x"F85C", x"F875",
    x"F88E", x"F8A7", x"F8C0", x"F8D9",
    x"F8F2", x"F90B", x"F924", x"F93D",
    x"F956", x"F96F", x"F988", x"F9A1",
    x"F9BA", x"F9D3", x"F9EC", x"FA05",
    x"FA1E", x"FA37", x"FA50", x"FA69",
    x"FA82", x"FA9B", x"FAB4", x"FACD",
    x"FAE6", x"FB00", x"FB19", x"FB32",
    x"FB4B", x"FB64", x"FB7D", x"FB96",
    x"FBAF", x"FBC8", x"FBE1", x"FBFA",
    x"FC13", x"FC2C", x"FC45", x"FC5F",
    x"FC78", x"FC91", x"FCAA", x"FCC3",
    x"FCDC", x"FCF5", x"FD0E", x"FD27",
    x"FD40", x"FD5A", x"FD73", x"FD8C",
    x"FDA5", x"FDBE", x"FDD7", x"FDF0",
    x"FE09", x"FE23", x"FE3C", x"FE55",
    x"FE6E", x"FE87", x"FEA0", x"FEB9",
    x"FED2", x"FEEC", x"FF05", x"FF1E",
    x"FF37", x"FF50", x"FF69", x"FF82",
    x"FF9B", x"FFB5", x"FFCE", x"FFE7");

signal angle, phase : signed(15 downto 0) := (others => '0');
signal turns, bin   : unsigned(15 downto 0) := (others => '0');
signal idx : integer  := 1; 

begin

angle <= signed(addr);
phase <= (angle + (shift_right(angle, 2) + shift_right(angle, 5) - shift_right(angle, 7)));
turns <= unsigned(phase); 
bin <= turns + to_unsigned(16, 16); 
idx <= to_integer( bin(15 downto 5));    

set_sine: process( idx ) 
begin 
  sine_out <= sine_table(idx);    
end process set_sine; 

end architecture behavioral; 
