library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; 
use work.array_types.all;

entity sine_lut is 
  port (
    clk_port : in std_logic; 
    cos_en   : in std_logic;  
    rads     : in std_logic_vector(15 downto 0); 
    sine     : out std_logic_vector(15 downto 0);
    set_port : out std_logic); -- 2.14 fixed point 
end entity sine_lut; 

architecture behavioral of sine_lut is 
  -- generate table from regfile decleration 
  constant sine_table : array_2048x16_t := (
    x"0000", x"0032", x"0065", x"0097",
    x"00C9", x"00FB", x"012E", x"0160",
    x"0192", x"01C4", x"01F7", x"0229",
    x"025B", x"028D", x"02C0", x"02F2",
    x"0324", x"0356", x"0388", x"03BB",
    x"03ED", x"041F", x"0451", x"0483",
    x"04B5", x"04E7", x"051A", x"054C",
    x"057E", x"05B0", x"05E2", x"0614",
    x"0646", x"0678", x"06AA", x"06DC",
    x"070E", x"0740", x"0772", x"07A4",
    x"07D6", x"0807", x"0839", x"086B",
    x"089D", x"08CF", x"0901", x"0932",
    x"0964", x"0996", x"09C7", x"09F9",
    x"0A2B", x"0A5C", x"0A8E", x"0AC0",
    x"0AF1", x"0B23", x"0B54", x"0B85",
    x"0BB7", x"0BE8", x"0C1A", x"0C4B",
    x"0C7C", x"0CAE", x"0CDF", x"0D10",
    x"0D41", x"0D72", x"0DA4", x"0DD5",
    x"0E06", x"0E37", x"0E68", x"0E99",
    x"0ECA", x"0EFB", x"0F2B", x"0F5C",
    x"0F8D", x"0FBE", x"0FEE", x"101F",
    x"1050", x"1080", x"10B1", x"10E1",
    x"1112", x"1142", x"1173", x"11A3",
    x"11D3", x"1204", x"1234", x"1264",
    x"1294", x"12C4", x"12F4", x"1324",
    x"1354", x"1384", x"13B4", x"13E4",
    x"1413", x"1443", x"1473", x"14A2",
    x"14D2", x"1501", x"1531", x"1560",
    x"1590", x"15BF", x"15EE", x"161D",
    x"164C", x"167C", x"16AB", x"16DA",
    x"1709", x"1737", x"1766", x"1795",
    x"17C4", x"17F2", x"1821", x"184F",
    x"187E", x"18AC", x"18DB", x"1909",
    x"1937", x"1965", x"1993", x"19C1",
    x"19EF", x"1A1D", x"1A4B", x"1A79",
    x"1AA7", x"1AD4", x"1B02", x"1B30",
    x"1B5D", x"1B8A", x"1BB8", x"1BE5",
    x"1C12", x"1C3F", x"1C6C", x"1C99",
    x"1CC6", x"1CF3", x"1D20", x"1D4D",
    x"1D79", x"1DA6", x"1DD3", x"1DFF",
    x"1E2B", x"1E58", x"1E84", x"1EB0",
    x"1EDC", x"1F08", x"1F34", x"1F60",
    x"1F8C", x"1FB7", x"1FE3", x"200F",
    x"203A", x"2065", x"2091", x"20BC",
    x"20E7", x"2112", x"213D", x"2168",
    x"2193", x"21BE", x"21E8", x"2213",
    x"223D", x"2268", x"2292", x"22BC",
    x"22E7", x"2311", x"233B", x"2365",
    x"238E", x"23B8", x"23E2", x"240B",
    x"2435", x"245E", x"2488", x"24B1",
    x"24DA", x"2503", x"252C", x"2555",
    x"257E", x"25A6", x"25CF", x"25F8",
    x"2620", x"2648", x"2671", x"2699",
    x"26C1", x"26E9", x"2711", x"2738",
    x"2760", x"2788", x"27AF", x"27D6",
    x"27FE", x"2825", x"284C", x"2873",
    x"289A", x"28C1", x"28E7", x"290E",
    x"2935", x"295B", x"2981", x"29A7",
    x"29CE", x"29F4", x"2A1A", x"2A3F",
    x"2A65", x"2A8B", x"2AB0", x"2AD6",
    x"2AFB", x"2B20", x"2B45", x"2B6A",
    x"2B8F", x"2BB4", x"2BD8", x"2BFD",
    x"2C21", x"2C46", x"2C6A", x"2C8E",
    x"2CB2", x"2CD6", x"2CFA", x"2D1E",
    x"2D41", x"2D65", x"2D88", x"2DAB",
    x"2DCF", x"2DF2", x"2E15", x"2E37",
    x"2E5A", x"2E7D", x"2E9F", x"2EC2",
    x"2EE4", x"2F06", x"2F28", x"2F4A",
    x"2F6C", x"2F8D", x"2FAF", x"2FD0",
    x"2FF2", x"3013", x"3034", x"3055",
    x"3076", x"3097", x"30B8", x"30D8",
    x"30F9", x"3119", x"3139", x"3159",
    x"3179", x"3199", x"31B9", x"31D8",
    x"31F8", x"3217", x"3236", x"3255",
    x"3274", x"3293", x"32B2", x"32D0",
    x"32EF", x"330D", x"332C", x"334A",
    x"3368", x"3386", x"33A3", x"33C1",
    x"33DF", x"33FC", x"3419", x"3436",
    x"3453", x"3470", x"348D", x"34AA",
    x"34C6", x"34E2", x"34FF", x"351B",
    x"3537", x"3553", x"356E", x"358A",
    x"35A5", x"35C1", x"35DC", x"35F7",
    x"3612", x"362D", x"3648", x"3662",
    x"367D", x"3697", x"36B1", x"36CB",
    x"36E5", x"36FF", x"3718", x"3732",
    x"374B", x"3765", x"377E", x"3797",
    x"37B0", x"37C8", x"37E1", x"37F9",
    x"3812", x"382A", x"3842", x"385A",
    x"3871", x"3889", x"38A1", x"38B8",
    x"38CF", x"38E6", x"38FD", x"3914",
    x"392B", x"3941", x"3958", x"396E",
    x"3984", x"399A", x"39B0", x"39C5",
    x"39DB", x"39F0", x"3A06", x"3A1B",
    x"3A30", x"3A45", x"3A59", x"3A6E",
    x"3A82", x"3A97", x"3AAB", x"3ABF",
    x"3AD3", x"3AE6", x"3AFA", x"3B0E",
    x"3B21", x"3B34", x"3B47", x"3B5A",
    x"3B6D", x"3B7F", x"3B92", x"3BA4",
    x"3BB6", x"3BC8", x"3BDA", x"3BEC",
    x"3BFD", x"3C0F", x"3C20", x"3C31",
    x"3C42", x"3C53", x"3C64", x"3C74",
    x"3C85", x"3C95", x"3CA5", x"3CB5",
    x"3CC5", x"3CD5", x"3CE4", x"3CF4",
    x"3D03", x"3D12", x"3D21", x"3D30",
    x"3D3F", x"3D4D", x"3D5B", x"3D6A",
    x"3D78", x"3D86", x"3D93", x"3DA1",
    x"3DAF", x"3DBC", x"3DC9", x"3DD6",
    x"3DE3", x"3DF0", x"3DFC", x"3E09",
    x"3E15", x"3E21", x"3E2D", x"3E39",
    x"3E45", x"3E50", x"3E5C", x"3E67",
    x"3E72", x"3E7D", x"3E88", x"3E92",
    x"3E9D", x"3EA7", x"3EB1", x"3EBB",
    x"3EC5", x"3ECF", x"3ED8", x"3EE2",
    x"3EEB", x"3EF4", x"3EFD", x"3F06",
    x"3F0F", x"3F17", x"3F20", x"3F28",
    x"3F30", x"3F38", x"3F40", x"3F47",
    x"3F4F", x"3F56", x"3F5D", x"3F64",
    x"3F6B", x"3F72", x"3F78", x"3F7F",
    x"3F85", x"3F8B", x"3F91", x"3F97",
    x"3F9C", x"3FA2", x"3FA7", x"3FAC",
    x"3FB1", x"3FB6", x"3FBB", x"3FBF",
    x"3FC4", x"3FC8", x"3FCC", x"3FD0",
    x"3FD4", x"3FD7", x"3FDB", x"3FDE",
    x"3FE1", x"3FE4", x"3FE7", x"3FEA",
    x"3FEC", x"3FEF", x"3FF1", x"3FF3",
    x"3FF5", x"3FF7", x"3FF8", x"3FFA",
    x"3FFB", x"3FFC", x"3FFD", x"3FFE",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFF", x"3FFF", x"3FFF",
    x"3FFF", x"3FFE", x"3FFD", x"3FFC",
    x"3FFB", x"3FFA", x"3FF8", x"3FF7",
    x"3FF5", x"3FF3", x"3FF1", x"3FEF",
    x"3FEC", x"3FEA", x"3FE7", x"3FE4",
    x"3FE1", x"3FDE", x"3FDB", x"3FD7",
    x"3FD4", x"3FD0", x"3FCC", x"3FC8",
    x"3FC4", x"3FBF", x"3FBB", x"3FB6",
    x"3FB1", x"3FAC", x"3FA7", x"3FA2",
    x"3F9C", x"3F97", x"3F91", x"3F8B",
    x"3F85", x"3F7F", x"3F78", x"3F72",
    x"3F6B", x"3F64", x"3F5D", x"3F56",
    x"3F4F", x"3F47", x"3F40", x"3F38",
    x"3F30", x"3F28", x"3F20", x"3F17",
    x"3F0F", x"3F06", x"3EFD", x"3EF4",
    x"3EEB", x"3EE2", x"3ED8", x"3ECF",
    x"3EC5", x"3EBB", x"3EB1", x"3EA7",
    x"3E9D", x"3E92", x"3E88", x"3E7D",
    x"3E72", x"3E67", x"3E5C", x"3E50",
    x"3E45", x"3E39", x"3E2D", x"3E21",
    x"3E15", x"3E09", x"3DFC", x"3DF0",
    x"3DE3", x"3DD6", x"3DC9", x"3DBC",
    x"3DAF", x"3DA1", x"3D93", x"3D86",
    x"3D78", x"3D6A", x"3D5B", x"3D4D",
    x"3D3F", x"3D30", x"3D21", x"3D12",
    x"3D03", x"3CF4", x"3CE4", x"3CD5",
    x"3CC5", x"3CB5", x"3CA5", x"3C95",
    x"3C85", x"3C74", x"3C64", x"3C53",
    x"3C42", x"3C31", x"3C20", x"3C0F",
    x"3BFD", x"3BEC", x"3BDA", x"3BC8",
    x"3BB6", x"3BA4", x"3B92", x"3B7F",
    x"3B6D", x"3B5A", x"3B47", x"3B34",
    x"3B21", x"3B0E", x"3AFA", x"3AE6",
    x"3AD3", x"3ABF", x"3AAB", x"3A97",
    x"3A82", x"3A6E", x"3A59", x"3A45",
    x"3A30", x"3A1B", x"3A06", x"39F0",
    x"39DB", x"39C5", x"39B0", x"399A",
    x"3984", x"396E", x"3958", x"3941",
    x"392B", x"3914", x"38FD", x"38E6",
    x"38CF", x"38B8", x"38A1", x"3889",
    x"3871", x"385A", x"3842", x"382A",
    x"3812", x"37F9", x"37E1", x"37C8",
    x"37B0", x"3797", x"377E", x"3765",
    x"374B", x"3732", x"3718", x"36FF",
    x"36E5", x"36CB", x"36B1", x"3697",
    x"367D", x"3662", x"3648", x"362D",
    x"3612", x"35F7", x"35DC", x"35C1",
    x"35A5", x"358A", x"356E", x"3553",
    x"3537", x"351B", x"34FF", x"34E2",
    x"34C6", x"34AA", x"348D", x"3470",
    x"3453", x"3436", x"3419", x"33FC",
    x"33DF", x"33C1", x"33A3", x"3386",
    x"3368", x"334A", x"332C", x"330D",
    x"32EF", x"32D0", x"32B2", x"3293",
    x"3274", x"3255", x"3236", x"3217",
    x"31F8", x"31D8", x"31B9", x"3199",
    x"3179", x"3159", x"3139", x"3119",
    x"30F9", x"30D8", x"30B8", x"3097",
    x"3076", x"3055", x"3034", x"3013",
    x"2FF2", x"2FD0", x"2FAF", x"2F8D",
    x"2F6C", x"2F4A", x"2F28", x"2F06",
    x"2EE4", x"2EC2", x"2E9F", x"2E7D",
    x"2E5A", x"2E37", x"2E15", x"2DF2",
    x"2DCF", x"2DAB", x"2D88", x"2D65",
    x"2D41", x"2D1E", x"2CFA", x"2CD6",
    x"2CB2", x"2C8E", x"2C6A", x"2C46",
    x"2C21", x"2BFD", x"2BD8", x"2BB4",
    x"2B8F", x"2B6A", x"2B45", x"2B20",
    x"2AFB", x"2AD6", x"2AB0", x"2A8B",
    x"2A65", x"2A3F", x"2A1A", x"29F4",
    x"29CE", x"29A7", x"2981", x"295B",
    x"2935", x"290E", x"28E7", x"28C1",
    x"289A", x"2873", x"284C", x"2825",
    x"27FE", x"27D6", x"27AF", x"2788",
    x"2760", x"2738", x"2711", x"26E9",
    x"26C1", x"2699", x"2671", x"2648",
    x"2620", x"25F8", x"25CF", x"25A6",
    x"257E", x"2555", x"252C", x"2503",
    x"24DA", x"24B1", x"2488", x"245E",
    x"2435", x"240B", x"23E2", x"23B8",
    x"238E", x"2365", x"233B", x"2311",
    x"22E7", x"22BC", x"2292", x"2268",
    x"223D", x"2213", x"21E8", x"21BE",
    x"2193", x"2168", x"213D", x"2112",
    x"20E7", x"20BC", x"2091", x"2065",
    x"203A", x"200F", x"1FE3", x"1FB7",
    x"1F8C", x"1F60", x"1F34", x"1F08",
    x"1EDC", x"1EB0", x"1E84", x"1E58",
    x"1E2B", x"1DFF", x"1DD3", x"1DA6",
    x"1D79", x"1D4D", x"1D20", x"1CF3",
    x"1CC6", x"1C99", x"1C6C", x"1C3F",
    x"1C12", x"1BE5", x"1BB8", x"1B8A",
    x"1B5D", x"1B30", x"1B02", x"1AD4",
    x"1AA7", x"1A79", x"1A4B", x"1A1D",
    x"19EF", x"19C1", x"1993", x"1965",
    x"1937", x"1909", x"18DB", x"18AC",
    x"187E", x"184F", x"1821", x"17F2",
    x"17C4", x"1795", x"1766", x"1737",
    x"1709", x"16DA", x"16AB", x"167C",
    x"164C", x"161D", x"15EE", x"15BF",
    x"1590", x"1560", x"1531", x"1501",
    x"14D2", x"14A2", x"1473", x"1443",
    x"1413", x"13E4", x"13B4", x"1384",
    x"1354", x"1324", x"12F4", x"12C4",
    x"1294", x"1264", x"1234", x"1204",
    x"11D3", x"11A3", x"1173", x"1142",
    x"1112", x"10E1", x"10B1", x"1080",
    x"1050", x"101F", x"0FEE", x"0FBE",
    x"0F8D", x"0F5C", x"0F2B", x"0EFB",
    x"0ECA", x"0E99", x"0E68", x"0E37",
    x"0E06", x"0DD5", x"0DA4", x"0D72",
    x"0D41", x"0D10", x"0CDF", x"0CAE",
    x"0C7C", x"0C4B", x"0C1A", x"0BE8",
    x"0BB7", x"0B85", x"0B54", x"0B23",
    x"0AF1", x"0AC0", x"0A8E", x"0A5C",
    x"0A2B", x"09F9", x"09C7", x"0996",
    x"0964", x"0932", x"0901", x"08CF",
    x"089D", x"086B", x"0839", x"0807",
    x"07D6", x"07A4", x"0772", x"0740",
    x"070E", x"06DC", x"06AA", x"0678",
    x"0646", x"0614", x"05E2", x"05B0",
    x"057E", x"054C", x"051A", x"04E7",
    x"04B5", x"0483", x"0451", x"041F",
    x"03ED", x"03BB", x"0388", x"0356",
    x"0324", x"02F2", x"02C0", x"028D",
    x"025B", x"0229", x"01F7", x"01C4",
    x"0192", x"0160", x"012E", x"00FB",
    x"00C9", x"0097", x"0065", x"0032",
    x"0000", x"FFCE", x"FF9B", x"FF69",
    x"FF37", x"FF05", x"FED2", x"FEA0",
    x"FE6E", x"FE3C", x"FE09", x"FDD7",
    x"FDA5", x"FD73", x"FD40", x"FD0E",
    x"FCDC", x"FCAA", x"FC78", x"FC45",
    x"FC13", x"FBE1", x"FBAF", x"FB7D",
    x"FB4B", x"FB19", x"FAE6", x"FAB4",
    x"FA82", x"FA50", x"FA1E", x"F9EC",
    x"F9BA", x"F988", x"F956", x"F924",
    x"F8F2", x"F8C0", x"F88E", x"F85C",
    x"F82A", x"F7F9", x"F7C7", x"F795",
    x"F763", x"F731", x"F6FF", x"F6CE",
    x"F69C", x"F66A", x"F639", x"F607",
    x"F5D5", x"F5A4", x"F572", x"F540",
    x"F50F", x"F4DD", x"F4AC", x"F47B",
    x"F449", x"F418", x"F3E6", x"F3B5",
    x"F384", x"F352", x"F321", x"F2F0",
    x"F2BF", x"F28E", x"F25C", x"F22B",
    x"F1FA", x"F1C9", x"F198", x"F167",
    x"F136", x"F105", x"F0D5", x"F0A4",
    x"F073", x"F042", x"F012", x"EFE1",
    x"EFB0", x"EF80", x"EF4F", x"EF1F",
    x"EEEE", x"EEBE", x"EE8D", x"EE5D",
    x"EE2D", x"EDFC", x"EDCC", x"ED9C",
    x"ED6C", x"ED3C", x"ED0C", x"ECDC",
    x"ECAC", x"EC7C", x"EC4C", x"EC1C",
    x"EBED", x"EBBD", x"EB8D", x"EB5E",
    x"EB2E", x"EAFF", x"EACF", x"EAA0",
    x"EA70", x"EA41", x"EA12", x"E9E3",
    x"E9B4", x"E984", x"E955", x"E926",
    x"E8F7", x"E8C9", x"E89A", x"E86B",
    x"E83C", x"E80E", x"E7DF", x"E7B1",
    x"E782", x"E754", x"E725", x"E6F7",
    x"E6C9", x"E69B", x"E66D", x"E63F",
    x"E611", x"E5E3", x"E5B5", x"E587",
    x"E559", x"E52C", x"E4FE", x"E4D0",
    x"E4A3", x"E476", x"E448", x"E41B",
    x"E3EE", x"E3C1", x"E394", x"E367",
    x"E33A", x"E30D", x"E2E0", x"E2B3",
    x"E287", x"E25A", x"E22D", x"E201",
    x"E1D5", x"E1A8", x"E17C", x"E150",
    x"E124", x"E0F8", x"E0CC", x"E0A0",
    x"E074", x"E049", x"E01D", x"DFF1",
    x"DFC6", x"DF9B", x"DF6F", x"DF44",
    x"DF19", x"DEEE", x"DEC3", x"DE98",
    x"DE6D", x"DE42", x"DE18", x"DDED",
    x"DDC3", x"DD98", x"DD6E", x"DD44",
    x"DD19", x"DCEF", x"DCC5", x"DC9B",
    x"DC72", x"DC48", x"DC1E", x"DBF5",
    x"DBCB", x"DBA2", x"DB78", x"DB4F",
    x"DB26", x"DAFD", x"DAD4", x"DAAB",
    x"DA82", x"DA5A", x"DA31", x"DA08",
    x"D9E0", x"D9B8", x"D98F", x"D967",
    x"D93F", x"D917", x"D8EF", x"D8C8",
    x"D8A0", x"D878", x"D851", x"D82A",
    x"D802", x"D7DB", x"D7B4", x"D78D",
    x"D766", x"D73F", x"D719", x"D6F2",
    x"D6CB", x"D6A5", x"D67F", x"D659",
    x"D632", x"D60C", x"D5E6", x"D5C1",
    x"D59B", x"D575", x"D550", x"D52A",
    x"D505", x"D4E0", x"D4BB", x"D496",
    x"D471", x"D44C", x"D428", x"D403",
    x"D3DF", x"D3BA", x"D396", x"D372",
    x"D34E", x"D32A", x"D306", x"D2E2",
    x"D2BF", x"D29B", x"D278", x"D255",
    x"D231", x"D20E", x"D1EB", x"D1C9",
    x"D1A6", x"D183", x"D161", x"D13E",
    x"D11C", x"D0FA", x"D0D8", x"D0B6",
    x"D094", x"D073", x"D051", x"D030",
    x"D00E", x"CFED", x"CFCC", x"CFAB",
    x"CF8A", x"CF69", x"CF48", x"CF28",
    x"CF07", x"CEE7", x"CEC7", x"CEA7",
    x"CE87", x"CE67", x"CE47", x"CE28",
    x"CE08", x"CDE9", x"CDCA", x"CDAB",
    x"CD8C", x"CD6D", x"CD4E", x"CD30",
    x"CD11", x"CCF3", x"CCD4", x"CCB6",
    x"CC98", x"CC7A", x"CC5D", x"CC3F",
    x"CC21", x"CC04", x"CBE7", x"CBCA",
    x"CBAD", x"CB90", x"CB73", x"CB56",
    x"CB3A", x"CB1E", x"CB01", x"CAE5",
    x"CAC9", x"CAAD", x"CA92", x"CA76",
    x"CA5B", x"CA3F", x"CA24", x"CA09",
    x"C9EE", x"C9D3", x"C9B8", x"C99E",
    x"C983", x"C969", x"C94F", x"C935",
    x"C91B", x"C901", x"C8E8", x"C8CE",
    x"C8B5", x"C89B", x"C882", x"C869",
    x"C850", x"C838", x"C81F", x"C807",
    x"C7EE", x"C7D6", x"C7BE", x"C7A6",
    x"C78F", x"C777", x"C75F", x"C748",
    x"C731", x"C71A", x"C703", x"C6EC",
    x"C6D5", x"C6BF", x"C6A8", x"C692",
    x"C67C", x"C666", x"C650", x"C63B",
    x"C625", x"C610", x"C5FA", x"C5E5",
    x"C5D0", x"C5BB", x"C5A7", x"C592",
    x"C57E", x"C569", x"C555", x"C541",
    x"C52D", x"C51A", x"C506", x"C4F2",
    x"C4DF", x"C4CC", x"C4B9", x"C4A6",
    x"C493", x"C481", x"C46E", x"C45C",
    x"C44A", x"C438", x"C426", x"C414",
    x"C403", x"C3F1", x"C3E0", x"C3CF",
    x"C3BE", x"C3AD", x"C39C", x"C38C",
    x"C37B", x"C36B", x"C35B", x"C34B",
    x"C33B", x"C32B", x"C31C", x"C30C",
    x"C2FD", x"C2EE", x"C2DF", x"C2D0",
    x"C2C1", x"C2B3", x"C2A5", x"C296",
    x"C288", x"C27A", x"C26D", x"C25F",
    x"C251", x"C244", x"C237", x"C22A",
    x"C21D", x"C210", x"C204", x"C1F7",
    x"C1EB", x"C1DF", x"C1D3", x"C1C7",
    x"C1BB", x"C1B0", x"C1A4", x"C199",
    x"C18E", x"C183", x"C178", x"C16E",
    x"C163", x"C159", x"C14F", x"C145",
    x"C13B", x"C131", x"C128", x"C11E",
    x"C115", x"C10C", x"C103", x"C0FA",
    x"C0F1", x"C0E9", x"C0E0", x"C0D8",
    x"C0D0", x"C0C8", x"C0C0", x"C0B9",
    x"C0B1", x"C0AA", x"C0A3", x"C09C",
    x"C095", x"C08E", x"C088", x"C081",
    x"C07B", x"C075", x"C06F", x"C069",
    x"C064", x"C05E", x"C059", x"C054",
    x"C04F", x"C04A", x"C045", x"C041",
    x"C03C", x"C038", x"C034", x"C030",
    x"C02C", x"C029", x"C025", x"C022",
    x"C01F", x"C01C", x"C019", x"C016",
    x"C014", x"C011", x"C00F", x"C00D",
    x"C00B", x"C009", x"C008", x"C006",
    x"C005", x"C004", x"C003", x"C002",
    x"C001", x"C001", x"C000", x"C000",
    x"C000", x"C000", x"C000", x"C001",
    x"C001", x"C002", x"C003", x"C004",
    x"C005", x"C006", x"C008", x"C009",
    x"C00B", x"C00D", x"C00F", x"C011",
    x"C014", x"C016", x"C019", x"C01C",
    x"C01F", x"C022", x"C025", x"C029",
    x"C02C", x"C030", x"C034", x"C038",
    x"C03C", x"C041", x"C045", x"C04A",
    x"C04F", x"C054", x"C059", x"C05E",
    x"C064", x"C069", x"C06F", x"C075",
    x"C07B", x"C081", x"C088", x"C08E",
    x"C095", x"C09C", x"C0A3", x"C0AA",
    x"C0B1", x"C0B9", x"C0C0", x"C0C8",
    x"C0D0", x"C0D8", x"C0E0", x"C0E9",
    x"C0F1", x"C0FA", x"C103", x"C10C",
    x"C115", x"C11E", x"C128", x"C131",
    x"C13B", x"C145", x"C14F", x"C159",
    x"C163", x"C16E", x"C178", x"C183",
    x"C18E", x"C199", x"C1A4", x"C1B0",
    x"C1BB", x"C1C7", x"C1D3", x"C1DF",
    x"C1EB", x"C1F7", x"C204", x"C210",
    x"C21D", x"C22A", x"C237", x"C244",
    x"C251", x"C25F", x"C26D", x"C27A",
    x"C288", x"C296", x"C2A5", x"C2B3",
    x"C2C1", x"C2D0", x"C2DF", x"C2EE",
    x"C2FD", x"C30C", x"C31C", x"C32B",
    x"C33B", x"C34B", x"C35B", x"C36B",
    x"C37B", x"C38C", x"C39C", x"C3AD",
    x"C3BE", x"C3CF", x"C3E0", x"C3F1",
    x"C403", x"C414", x"C426", x"C438",
    x"C44A", x"C45C", x"C46E", x"C481",
    x"C493", x"C4A6", x"C4B9", x"C4CC",
    x"C4DF", x"C4F2", x"C506", x"C51A",
    x"C52D", x"C541", x"C555", x"C569",
    x"C57E", x"C592", x"C5A7", x"C5BB",
    x"C5D0", x"C5E5", x"C5FA", x"C610",
    x"C625", x"C63B", x"C650", x"C666",
    x"C67C", x"C692", x"C6A8", x"C6BF",
    x"C6D5", x"C6EC", x"C703", x"C71A",
    x"C731", x"C748", x"C75F", x"C777",
    x"C78F", x"C7A6", x"C7BE", x"C7D6",
    x"C7EE", x"C807", x"C81F", x"C838",
    x"C850", x"C869", x"C882", x"C89B",
    x"C8B5", x"C8CE", x"C8E8", x"C901",
    x"C91B", x"C935", x"C94F", x"C969",
    x"C983", x"C99E", x"C9B8", x"C9D3",
    x"C9EE", x"CA09", x"CA24", x"CA3F",
    x"CA5B", x"CA76", x"CA92", x"CAAD",
    x"CAC9", x"CAE5", x"CB01", x"CB1E",
    x"CB3A", x"CB56", x"CB73", x"CB90",
    x"CBAD", x"CBCA", x"CBE7", x"CC04",
    x"CC21", x"CC3F", x"CC5D", x"CC7A",
    x"CC98", x"CCB6", x"CCD4", x"CCF3",
    x"CD11", x"CD30", x"CD4E", x"CD6D",
    x"CD8C", x"CDAB", x"CDCA", x"CDE9",
    x"CE08", x"CE28", x"CE47", x"CE67",
    x"CE87", x"CEA7", x"CEC7", x"CEE7",
    x"CF07", x"CF28", x"CF48", x"CF69",
    x"CF8A", x"CFAB", x"CFCC", x"CFED",
    x"D00E", x"D030", x"D051", x"D073",
    x"D094", x"D0B6", x"D0D8", x"D0FA",
    x"D11C", x"D13E", x"D161", x"D183",
    x"D1A6", x"D1C9", x"D1EB", x"D20E",
    x"D231", x"D255", x"D278", x"D29B",
    x"D2BF", x"D2E2", x"D306", x"D32A",
    x"D34E", x"D372", x"D396", x"D3BA",
    x"D3DF", x"D403", x"D428", x"D44C",
    x"D471", x"D496", x"D4BB", x"D4E0",
    x"D505", x"D52A", x"D550", x"D575",
    x"D59B", x"D5C1", x"D5E6", x"D60C",
    x"D632", x"D659", x"D67F", x"D6A5",
    x"D6CB", x"D6F2", x"D719", x"D73F",
    x"D766", x"D78D", x"D7B4", x"D7DB",
    x"D802", x"D82A", x"D851", x"D878",
    x"D8A0", x"D8C8", x"D8EF", x"D917",
    x"D93F", x"D967", x"D98F", x"D9B8",
    x"D9E0", x"DA08", x"DA31", x"DA5A",
    x"DA82", x"DAAB", x"DAD4", x"DAFD",
    x"DB26", x"DB4F", x"DB78", x"DBA2",
    x"DBCB", x"DBF5", x"DC1E", x"DC48",
    x"DC72", x"DC9B", x"DCC5", x"DCEF",
    x"DD19", x"DD44", x"DD6E", x"DD98",
    x"DDC3", x"DDED", x"DE18", x"DE42",
    x"DE6D", x"DE98", x"DEC3", x"DEEE",
    x"DF19", x"DF44", x"DF6F", x"DF9B",
    x"DFC6", x"DFF1", x"E01D", x"E049",
    x"E074", x"E0A0", x"E0CC", x"E0F8",
    x"E124", x"E150", x"E17C", x"E1A8",
    x"E1D5", x"E201", x"E22D", x"E25A",
    x"E287", x"E2B3", x"E2E0", x"E30D",
    x"E33A", x"E367", x"E394", x"E3C1",
    x"E3EE", x"E41B", x"E448", x"E476",
    x"E4A3", x"E4D0", x"E4FE", x"E52C",
    x"E559", x"E587", x"E5B5", x"E5E3",
    x"E611", x"E63F", x"E66D", x"E69B",
    x"E6C9", x"E6F7", x"E725", x"E754",
    x"E782", x"E7B1", x"E7DF", x"E80E",
    x"E83C", x"E86B", x"E89A", x"E8C9",
    x"E8F7", x"E926", x"E955", x"E984",
    x"E9B4", x"E9E3", x"EA12", x"EA41",
    x"EA70", x"EAA0", x"EACF", x"EAFF",
    x"EB2E", x"EB5E", x"EB8D", x"EBBD",
    x"EBED", x"EC1C", x"EC4C", x"EC7C",
    x"ECAC", x"ECDC", x"ED0C", x"ED3C",
    x"ED6C", x"ED9C", x"EDCC", x"EDFC",
    x"EE2D", x"EE5D", x"EE8D", x"EEBE",
    x"EEEE", x"EF1F", x"EF4F", x"EF80",
    x"EFB0", x"EFE1", x"F012", x"F042",
    x"F073", x"F0A4", x"F0D5", x"F105",
    x"F136", x"F167", x"F198", x"F1C9",
    x"F1FA", x"F22B", x"F25C", x"F28E",
    x"F2BF", x"F2F0", x"F321", x"F352",
    x"F384", x"F3B5", x"F3E6", x"F418",
    x"F449", x"F47B", x"F4AC", x"F4DD",
    x"F50F", x"F540", x"F572", x"F5A4",
    x"F5D5", x"F607", x"F639", x"F66A",
    x"F69C", x"F6CE", x"F6FF", x"F731",
    x"F763", x"F795", x"F7C7", x"F7F9",
    x"F82A", x"F85C", x"F88E", x"F8C0",
    x"F8F2", x"F924", x"F956", x"F988",
    x"F9BA", x"F9EC", x"FA1E", x"FA50",
    x"FA82", x"FAB4", x"FAE6", x"FB19",
    x"FB4B", x"FB7D", x"FBAF", x"FBE1",
    x"FC13", x"FC45", x"FC78", x"FCAA",
    x"FCDC", x"FD0E", x"FD40", x"FD73",
    x"FDA5", x"FDD7", x"FE09", x"FE3C",
    x"FE6E", x"FEA0", x"FED2", x"FF05",
    x"FF37", x"FF69", x"FF9B", x"FFCE");

signal angle, phase : signed(15 downto 0)   := (others => '0');
signal turns, bin   : unsigned(15 downto 0) := (others => '0');
signal idx          : integer := 1; 

begin

angle <= signed(rads);
phase <= shift_left((angle + (shift_right(angle, 2) + shift_right(angle, 5) - shift_right(angle, 7))), 1);

-- handle cosine internally by adding turns to phase (specific to 2048 value table)  
turns <=  unsigned(phase)          when cos_en = '1' else  
         (unsigned(phase) + 16384) when cos_en = '0'; 
bin   <= turns + 16; 
idx   <= to_integer( bin(15 downto 5));    

-- set read value on ff and assert that value can be read
set_sine: process( clk_port ) 
begin 
  if rising_edge( clk_port ) then
    set_port <= '1';
    sine     <= sine_table(idx);    
  end if; 
end process set_sine; 

end architecture behavioral; 
