library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; 
use work.array_types.all;

entity newton_lut is 
  port (
    clk_port : in std_logic; 
    addr     : in std_logic_vector(9 downto 0); 
    seed     : out std_logic_vector(23 downto 0); -- 6.17 signed fixed point 
    set_port : out std_logic);  
end entity newton_lut; 

architecture behavioral of newton_lut is 
  constant newton_table : array_1024x24_t := ( 
    x"01FFC0", x"01FF40", x"01FEC1", x"01FE42",
    x"01FDC3", x"01FD44", x"01FCC5", x"01FC47",
    x"01FBC9", x"01FB4B", x"01FACE", x"01FA50",
    x"01F9D3", x"01F956", x"01F8DA", x"01F85E",
    x"01F7E1", x"01F766", x"01F6EA", x"01F66F",
    x"01F5F4", x"01F579", x"01F4FE", x"01F483",
    x"01F409", x"01F38F", x"01F316", x"01F29C",
    x"01F223", x"01F1AA", x"01F131", x"01F0B8",
    x"01F040", x"01EFC8", x"01EF50", x"01EED8",
    x"01EE61", x"01EDEA", x"01ED73", x"01ECFC",
    x"01EC85", x"01EC0F", x"01EB99", x"01EB23",
    x"01EAAD", x"01EA38", x"01E9C3", x"01E94E",
    x"01E8D9", x"01E864", x"01E7F0", x"01E77C",
    x"01E708", x"01E694", x"01E621", x"01E5AD",
    x"01E53A", x"01E4C7", x"01E455", x"01E3E2",
    x"01E370", x"01E2FE", x"01E28C", x"01E21B",
    x"01E1A9", x"01E138", x"01E0C7", x"01E056",
    x"01DFE6", x"01DF75", x"01DF05", x"01DE95",
    x"01DE26", x"01DDB6", x"01DD47", x"01DCD8",
    x"01DC69", x"01DBFA", x"01DB8B", x"01DB1D",
    x"01DAAF", x"01DA41", x"01D9D3", x"01D966",
    x"01D8F8", x"01D88B", x"01D81E", x"01D7B2",
    x"01D745", x"01D6D9", x"01D66D", x"01D601",
    x"01D595", x"01D529", x"01D4BE", x"01D453",
    x"01D3E8", x"01D37D", x"01D312", x"01D2A8",
    x"01D23E", x"01D1D4", x"01D16A", x"01D100",
    x"01D097", x"01D02D", x"01CFC4", x"01CF5B",
    x"01CEF3", x"01CE8A", x"01CE22", x"01CDB9",
    x"01CD51", x"01CCEA", x"01CC82", x"01CC1B",
    x"01CBB3", x"01CB4C", x"01CAE5", x"01CA7E",
    x"01CA18", x"01C9B2", x"01C94B", x"01C8E5",
    x"01C87F", x"01C81A", x"01C7B4", x"01C74F",
    x"01C6EA", x"01C685", x"01C620", x"01C5BC",
    x"01C557", x"01C4F3", x"01C48F", x"01C42B",
    x"01C3C7", x"01C364", x"01C300", x"01C29D",
    x"01C23A", x"01C1D7", x"01C174", x"01C112",
    x"01C0AF", x"01C04D", x"01BFEB", x"01BF89",
    x"01BF27", x"01BEC6", x"01BE64", x"01BE03",
    x"01BDA2", x"01BD41", x"01BCE1", x"01BC80",
    x"01BC20", x"01BBBF", x"01BB5F", x"01BAFF",
    x"01BAA0", x"01BA40", x"01B9E1", x"01B981",
    x"01B922", x"01B8C3", x"01B865", x"01B806",
    x"01B7A8", x"01B749", x"01B6EB", x"01B68D",
    x"01B62F", x"01B5D2", x"01B574", x"01B517",
    x"01B4BA", x"01B45C", x"01B400", x"01B3A3",
    x"01B346", x"01B2EA", x"01B28E", x"01B231",
    x"01B1D5", x"01B17A", x"01B11E", x"01B0C2",
    x"01B067", x"01B00C", x"01AFB1", x"01AF56",
    x"01AEFB", x"01AEA0", x"01AE46", x"01ADEC",
    x"01AD91", x"01AD37", x"01ACDE", x"01AC84",
    x"01AC2A", x"01ABD1", x"01AB77", x"01AB1E",
    x"01AAC5", x"01AA6C", x"01AA14", x"01A9BB",
    x"01A963", x"01A90A", x"01A8B2", x"01A85A",
    x"01A802", x"01A7AB", x"01A753", x"01A6FC",
    x"01A6A4", x"01A64D", x"01A5F6", x"01A59F",
    x"01A549", x"01A4F2", x"01A49C", x"01A445",
    x"01A3EF", x"01A399", x"01A343", x"01A2ED",
    x"01A298", x"01A242", x"01A1ED", x"01A198",
    x"01A143", x"01A0EE", x"01A099", x"01A044",
    x"019FF0", x"019F9B", x"019F47", x"019EF3",
    x"019E9F", x"019E4B", x"019DF7", x"019DA4",
    x"019D50", x"019CFD", x"019CAA", x"019C57",
    x"019C04", x"019BB1", x"019B5E", x"019B0C",
    x"019AB9", x"019A67", x"019A15", x"0199C3",
    x"019971", x"01991F", x"0198CD", x"01987C",
    x"01982A", x"0197D9", x"019788", x"019737",
    x"0196E6", x"019695", x"019644", x"0195F4",
    x"0195A4", x"019553", x"019503", x"0194B3",
    x"019463", x"019413", x"0193C4", x"019374",
    x"019325", x"0192D5", x"019286", x"019237",
    x"0191E8", x"019199", x"01914B", x"0190FC",
    x"0190AE", x"01905F", x"019011", x"018FC3",
    x"018F75", x"018F27", x"018EDA", x"018E8C",
    x"018E3E", x"018DF1", x"018DA4", x"018D57",
    x"018D0A", x"018CBD", x"018C70", x"018C23",
    x"018BD7", x"018B8A", x"018B3E", x"018AF2",
    x"018AA6", x"018A5A", x"018A0E", x"0189C2",
    x"018976", x"01892B", x"0188DF", x"018894",
    x"018849", x"0187FE", x"0187B3", x"018768",
    x"01871D", x"0186D2", x"018688", x"01863E",
    x"0185F3", x"0185A9", x"01855F", x"018515",
    x"0184CB", x"018481", x"018438", x"0183EE",
    x"0183A5", x"01835B", x"018312", x"0182C9",
    x"018280", x"018237", x"0181EE", x"0181A6",
    x"01815D", x"018115", x"0180CC", x"018084",
    x"01803C", x"017FF4", x"017FAC", x"017F64",
    x"017F1D", x"017ED5", x"017E8D", x"017E46",
    x"017DFF", x"017DB7", x"017D70", x"017D29",
    x"017CE3", x"017C9C", x"017C55", x"017C0E",
    x"017BC8", x"017B82", x"017B3B", x"017AF5",
    x"017AAF", x"017A69", x"017A23", x"0179DD",
    x"017998", x"017952", x"01790D", x"0178C7",
    x"017882", x"01783D", x"0177F8", x"0177B3",
    x"01776E", x"017729", x"0176E5", x"0176A0",
    x"01765C", x"017617", x"0175D3", x"01758F",
    x"01754B", x"017507", x"0174C3", x"01747F",
    x"01743B", x"0173F8", x"0173B4", x"017371",
    x"01732D", x"0172EA", x"0172A7", x"017264",
    x"017221", x"0171DE", x"01719B", x"017159",
    x"017116", x"0170D4", x"017091", x"01704F",
    x"01700D", x"016FCB", x"016F89", x"016F47",
    x"016F05", x"016EC3", x"016E82", x"016E40",
    x"016DFF", x"016DBD", x"016D7C", x"016D3B",
    x"016CFA", x"016CB9", x"016C78", x"016C37",
    x"016BF6", x"016BB6", x"016B75", x"016B35",
    x"016AF4", x"016AB4", x"016A74", x"016A34",
    x"0169F4", x"0169B4", x"016974", x"016934",
    x"0168F5", x"0168B5", x"016876", x"016836",
    x"0167F7", x"0167B8", x"016778", x"016739",
    x"0166FA", x"0166BC", x"01667D", x"01663E",
    x"0165FF", x"0165C1", x"016582", x"016544",
    x"016506", x"0164C8", x"01648A", x"01644C",
    x"01640E", x"0163D0", x"016392", x"016354",
    x"016317", x"0162D9", x"01629C", x"01625E",
    x"016221", x"0161E4", x"0161A7", x"01616A",
    x"01612D", x"0160F0", x"0160B3", x"016076",
    x"01603A", x"015FFD", x"015FC1", x"015F84",
    x"015F48", x"015F0C", x"015ED0", x"015E94",
    x"015E58", x"015E1C", x"015DE0", x"015DA4",
    x"015D69", x"015D2D", x"015CF2", x"015CB6",
    x"015C7B", x"015C40", x"015C04", x"015BC9",
    x"015B8E", x"015B53", x"015B18", x"015ADE",
    x"015AA3", x"015A68", x"015A2E", x"0159F3",
    x"0159B9", x"01597F", x"015944", x"01590A",
    x"0158D0", x"015896", x"01585C", x"015822",
    x"0157E8", x"0157AF", x"015775", x"01573C",
    x"015702", x"0156C9", x"01568F", x"015656",
    x"01561D", x"0155E4", x"0155AB", x"015572",
    x"015539", x"015500", x"0154C7", x"01548F",
    x"015456", x"01541E", x"0153E5", x"0153AD",
    x"015374", x"01533C", x"015304", x"0152CC",
    x"015294", x"01525C", x"015224", x"0151EC",
    x"0151B5", x"01517D", x"015145", x"01510E",
    x"0150D6", x"01509F", x"015068", x"015031",
    x"014FF9", x"014FC2", x"014F8B", x"014F54",
    x"014F1E", x"014EE7", x"014EB0", x"014E79",
    x"014E43", x"014E0C", x"014DD6", x"014D9F",
    x"014D69", x"014D33", x"014CFD", x"014CC7",
    x"014C91", x"014C5B", x"014C25", x"014BEF",
    x"014BB9", x"014B83", x"014B4E", x"014B18",
    x"014AE3", x"014AAD", x"014A78", x"014A43",
    x"014A0D", x"0149D8", x"0149A3", x"01496E",
    x"014939", x"014904", x"0148CF", x"01489B",
    x"014866", x"014831", x"0147FD", x"0147C8",
    x"014794", x"014760", x"01472B", x"0146F7",
    x"0146C3", x"01468F", x"01465B", x"014627",
    x"0145F3", x"0145BF", x"01458B", x"014557",
    x"014524", x"0144F0", x"0144BD", x"014489",
    x"014456", x"014423", x"0143EF", x"0143BC",
    x"014389", x"014356", x"014323", x"0142F0",
    x"0142BD", x"01428A", x"014257", x"014225",
    x"0141F2", x"0141BF", x"01418D", x"01415A",
    x"014128", x"0140F6", x"0140C3", x"014091",
    x"01405F", x"01402D", x"013FFB", x"013FC9",
    x"013F97", x"013F65", x"013F34", x"013F02",
    x"013ED0", x"013E9F", x"013E6D", x"013E3C",
    x"013E0A", x"013DD9", x"013DA7", x"013D76",
    x"013D45", x"013D14", x"013CE3", x"013CB2",
    x"013C81", x"013C50", x"013C1F", x"013BEE",
    x"013BBE", x"013B8D", x"013B5C", x"013B2C",
    x"013AFB", x"013ACB", x"013A9B", x"013A6A",
    x"013A3A", x"013A0A", x"0139DA", x"0139AA",
    x"01397A", x"01394A", x"01391A", x"0138EA",
    x"0138BA", x"01388B", x"01385B", x"01382B",
    x"0137FC", x"0137CC", x"01379D", x"01376D",
    x"01373E", x"01370F", x"0136E0", x"0136B0",
    x"013681", x"013652", x"013623", x"0135F4",
    x"0135C5", x"013597", x"013568", x"013539",
    x"01350A", x"0134DC", x"0134AD", x"01347F",
    x"013450", x"013422", x"0133F4", x"0133C5",
    x"013397", x"013369", x"01333B", x"01330D",
    x"0132DF", x"0132B1", x"013283", x"013255",
    x"013227", x"0131FA", x"0131CC", x"01319E",
    x"013171", x"013143", x"013116", x"0130E8",
    x"0130BB", x"01308E", x"013060", x"013033",
    x"013006", x"012FD9", x"012FAC", x"012F7F",
    x"012F52", x"012F25", x"012EF8", x"012ECB",
    x"012E9F", x"012E72", x"012E45", x"012E19",
    x"012DEC", x"012DC0", x"012D93", x"012D67",
    x"012D3A", x"012D0E", x"012CE2", x"012CB6",
    x"012C8A", x"012C5E", x"012C32", x"012C06",
    x"012BDA", x"012BAE", x"012B82", x"012B56",
    x"012B2A", x"012AFF", x"012AD3", x"012AA8",
    x"012A7C", x"012A51", x"012A25", x"0129FA",
    x"0129CE", x"0129A3", x"012978", x"01294D",
    x"012922", x"0128F7", x"0128CB", x"0128A0",
    x"012876", x"01284B", x"012820", x"0127F5",
    x"0127CA", x"0127A0", x"012775", x"01274A",
    x"012720", x"0126F5", x"0126CB", x"0126A0",
    x"012676", x"01264C", x"012621", x"0125F7",
    x"0125CD", x"0125A3", x"012579", x"01254F",
    x"012525", x"0124FB", x"0124D1", x"0124A7",
    x"01247D", x"012454", x"01242A", x"012400",
    x"0123D7", x"0123AD", x"012384", x"01235A",
    x"012331", x"012307", x"0122DE", x"0122B5",
    x"01228B", x"012262", x"012239", x"012210",
    x"0121E7", x"0121BE", x"012195", x"01216C",
    x"012143", x"01211A", x"0120F2", x"0120C9",
    x"0120A0", x"012077", x"01204F", x"012026",
    x"011FFE", x"011FD5", x"011FAD", x"011F84",
    x"011F5C", x"011F34", x"011F0C", x"011EE3",
    x"011EBB", x"011E93", x"011E6B", x"011E43",
    x"011E1B", x"011DF3", x"011DCB", x"011DA3",
    x"011D7B", x"011D54", x"011D2C", x"011D04",
    x"011CDD", x"011CB5", x"011C8D", x"011C66",
    x"011C3E", x"011C17", x"011BF0", x"011BC8",
    x"011BA1", x"011B7A", x"011B53", x"011B2B",
    x"011B04", x"011ADD", x"011AB6", x"011A8F",
    x"011A68", x"011A41", x"011A1A", x"0119F3",
    x"0119CD", x"0119A6", x"01197F", x"011959",
    x"011932", x"01190B", x"0118E5", x"0118BE",
    x"011898", x"011871", x"01184B", x"011825",
    x"0117FE", x"0117D8", x"0117B2", x"01178C",
    x"011766", x"01173F", x"011719", x"0116F3",
    x"0116CD", x"0116A7", x"011682", x"01165C",
    x"011636", x"011610", x"0115EA", x"0115C5",
    x"01159F", x"011579", x"011554", x"01152E",
    x"011509", x"0114E3", x"0114BE", x"011499",
    x"011473", x"01144E", x"011429", x"011404",
    x"0113DE", x"0113B9", x"011394", x"01136F",
    x"01134A", x"011325", x"011300", x"0112DB",
    x"0112B6", x"011291", x"01126D", x"011248",
    x"011223", x"0111FF", x"0111DA", x"0111B5",
    x"011191", x"01116C", x"011148", x"011123",
    x"0110FF", x"0110DA", x"0110B6", x"011092",
    x"01106E", x"011049", x"011025", x"011001",
    x"010FDD", x"010FB9", x"010F95", x"010F71",
    x"010F4D", x"010F29", x"010F05", x"010EE1",
    x"010EBD", x"010E9A", x"010E76", x"010E52",
    x"010E2F", x"010E0B", x"010DE7", x"010DC4",
    x"010DA0", x"010D7D", x"010D59", x"010D36",
    x"010D13", x"010CEF", x"010CCC", x"010CA9",
    x"010C85", x"010C62", x"010C3F", x"010C1C",
    x"010BF9", x"010BD6", x"010BB3", x"010B90",
    x"010B6D", x"010B4A", x"010B27", x"010B04",
    x"010AE2", x"010ABF", x"010A9C", x"010A79",
    x"010A57", x"010A34", x"010A12", x"0109EF",
    x"0109CC", x"0109AA", x"010988", x"010965",
    x"010943", x"010920", x"0108FE", x"0108DC",
    x"0108BA", x"010897", x"010875", x"010853",
    x"010831", x"01080F", x"0107ED", x"0107CB",
    x"0107A9", x"010787", x"010765", x"010743",
    x"010721", x"010700", x"0106DE", x"0106BC",
    x"01069B", x"010679", x"010657", x"010636",
    x"010614", x"0105F3", x"0105D1", x"0105B0",
    x"01058E", x"01056D", x"01054B", x"01052A",
    x"010509", x"0104E8", x"0104C6", x"0104A5",
    x"010484", x"010463", x"010442", x"010421",
    x"010400", x"0103DF", x"0103BE", x"01039D",
    x"01037C", x"01035B", x"01033A", x"010319",
    x"0102F9", x"0102D8", x"0102B7", x"010297",
    x"010276", x"010255", x"010235", x"010214",
    x"0101F4", x"0101D3", x"0101B3", x"010192",
    x"010172", x"010152", x"010131", x"010111",
    x"0100F1", x"0100D1", x"0100B0", x"010090",
    x"010070", x"010050", x"010030", x"010010"
  );
  signal uAddr : unsigned(9 downto 0) := (others => '0'); 
  signal idx   : integer := 0; 
begin 

-- get integer index 
uAddr <= unsigned(addr);
idx   <= to_integer(uAddr);

-- set read value in flop 
set_seed: process( clk_port )
begin 
  if rising_edge( clk_port ) then 
    set_port <= '1'; 
    seed     <= newton_table(idx);
  end if; 
end process set_seed; 

end architecture behavioral;
